
module weights_rom_depthwise_pointwise_3 (
    input wire [15:0] addr, 
    output reg [7:0] data) ;
    reg [7:0] rom [0:36863] ; 
    initial
        begin
            rom[0] = 8'he3 ;
            rom[1] = 8'hec ;
            rom[2] = 8'h2b ;
            rom[3] = 8'he0 ;
            rom[4] = 8'h05 ;
            rom[5] = 8'h09 ;
            rom[6] = 8'h10 ;
            rom[7] = 8'h04 ;
            rom[8] = 8'he6 ;
            rom[9] = 8'h0b ;
            rom[10] = 8'he3 ;
            rom[11] = 8'hdb ;
            rom[12] = 8'h0f ;
            rom[13] = 8'hfd ;
            rom[14] = 8'h18 ;
            rom[15] = 8'hde ;
            rom[16] = 8'h19 ;
            rom[17] = 8'hdb ;
            rom[18] = 8'he5 ;
            rom[19] = 8'hf2 ;
            rom[20] = 8'h20 ;
            rom[21] = 8'hfd ;
            rom[22] = 8'h1a ;
            rom[23] = 8'he1 ;
            rom[24] = 8'hf7 ;
            rom[25] = 8'hfa ;
            rom[26] = 8'h02 ;
            rom[27] = 8'hf9 ;
            rom[28] = 8'h01 ;
            rom[29] = 8'hf6 ;
            rom[30] = 8'h02 ;
            rom[31] = 8'h0f ;
            rom[32] = 8'hf9 ;
            rom[33] = 8'h03 ;
            rom[34] = 8'hea ;
            rom[35] = 8'hd7 ;
            rom[36] = 8'h22 ;
            rom[37] = 8'h06 ;
            rom[38] = 8'h01 ;
            rom[39] = 8'h02 ;
            rom[40] = 8'hff ;
            rom[41] = 8'hf0 ;
            rom[42] = 8'h19 ;
            rom[43] = 8'hda ;
            rom[44] = 8'h1f ;
            rom[45] = 8'h0b ;
            rom[46] = 8'h05 ;
            rom[47] = 8'hee ;
            rom[48] = 8'h1f ;
            rom[49] = 8'h0c ;
            rom[50] = 8'hdc ;
            rom[51] = 8'hf8 ;
            rom[52] = 8'hfa ;
            rom[53] = 8'hf2 ;
            rom[54] = 8'hcc ;
            rom[55] = 8'hd9 ;
            rom[56] = 8'h0e ;
            rom[57] = 8'h0b ;
            rom[58] = 8'h05 ;
            rom[59] = 8'h21 ;
            rom[60] = 8'h12 ;
            rom[61] = 8'hd9 ;
            rom[62] = 8'hda ;
            rom[63] = 8'he4 ;
            rom[64] = 8'h09 ;
            rom[65] = 8'h0a ;
            rom[66] = 8'h1e ;
            rom[67] = 8'he2 ;
            rom[68] = 8'hd4 ;
            rom[69] = 8'hee ;
            rom[70] = 8'hfb ;
            rom[71] = 8'he2 ;
            rom[72] = 8'h18 ;
            rom[73] = 8'hf2 ;
            rom[74] = 8'hcf ;
            rom[75] = 8'h1b ;
            rom[76] = 8'hf4 ;
            rom[77] = 8'h04 ;
            rom[78] = 8'he5 ;
            rom[79] = 8'h26 ;
            rom[80] = 8'h0b ;
            rom[81] = 8'h27 ;
            rom[82] = 8'hdb ;
            rom[83] = 8'h06 ;
            rom[84] = 8'hf6 ;
            rom[85] = 8'h0b ;
            rom[86] = 8'h15 ;
            rom[87] = 8'hc5 ;
            rom[88] = 8'hf9 ;
            rom[89] = 8'he9 ;
            rom[90] = 8'h0a ;
            rom[91] = 8'h05 ;
            rom[92] = 8'hff ;
            rom[93] = 8'h15 ;
            rom[94] = 8'hdd ;
            rom[95] = 8'hf1 ;
            rom[96] = 8'hfb ;
            rom[97] = 8'hfb ;
            rom[98] = 8'hd7 ;
            rom[99] = 8'h0e ;
            rom[100] = 8'h1a ;
            rom[101] = 8'he7 ;
            rom[102] = 8'hf3 ;
            rom[103] = 8'hf1 ;
            rom[104] = 8'he1 ;
            rom[105] = 8'h01 ;
            rom[106] = 8'hfc ;
            rom[107] = 8'hfa ;
            rom[108] = 8'h10 ;
            rom[109] = 8'hee ;
            rom[110] = 8'h24 ;
            rom[111] = 8'hd7 ;
            rom[112] = 8'hef ;
            rom[113] = 8'h0d ;
            rom[114] = 8'he6 ;
            rom[115] = 8'hda ;
            rom[116] = 8'h25 ;
            rom[117] = 8'hd6 ;
            rom[118] = 8'h11 ;
            rom[119] = 8'h00 ;
            rom[120] = 8'hce ;
            rom[121] = 8'hf7 ;
            rom[122] = 8'h1f ;
            rom[123] = 8'hf1 ;
            rom[124] = 8'hdc ;
            rom[125] = 8'hd5 ;
            rom[126] = 8'hcf ;
            rom[127] = 8'hea ;
            rom[128] = 8'h13 ;
            rom[129] = 8'h10 ;
            rom[130] = 8'h0f ;
            rom[131] = 8'h07 ;
            rom[132] = 8'h06 ;
            rom[133] = 8'he5 ;
            rom[134] = 8'h0a ;
            rom[135] = 8'hf0 ;
            rom[136] = 8'h02 ;
            rom[137] = 8'hf9 ;
            rom[138] = 8'h09 ;
            rom[139] = 8'h1c ;
            rom[140] = 8'h1c ;
            rom[141] = 8'h12 ;
            rom[142] = 8'hdb ;
            rom[143] = 8'h12 ;
            rom[144] = 8'he3 ;
            rom[145] = 8'hef ;
            rom[146] = 8'he7 ;
            rom[147] = 8'he8 ;
            rom[148] = 8'he7 ;
            rom[149] = 8'hef ;
            rom[150] = 8'hce ;
            rom[151] = 8'hda ;
            rom[152] = 8'he2 ;
            rom[153] = 8'h15 ;
            rom[154] = 8'hf0 ;
            rom[155] = 8'hbb ;
            rom[156] = 8'h1c ;
            rom[157] = 8'hca ;
            rom[158] = 8'hdb ;
            rom[159] = 8'he2 ;
            rom[160] = 8'hd8 ;
            rom[161] = 8'hf5 ;
            rom[162] = 8'hf0 ;
            rom[163] = 8'h1f ;
            rom[164] = 8'hd3 ;
            rom[165] = 8'hed ;
            rom[166] = 8'he2 ;
            rom[167] = 8'he3 ;
            rom[168] = 8'hfa ;
            rom[169] = 8'hfc ;
            rom[170] = 8'h1e ;
            rom[171] = 8'hbf ;
            rom[172] = 8'hf8 ;
            rom[173] = 8'he7 ;
            rom[174] = 8'hf6 ;
            rom[175] = 8'hf6 ;
            rom[176] = 8'hd4 ;
            rom[177] = 8'he0 ;
            rom[178] = 8'hdf ;
            rom[179] = 8'h04 ;
            rom[180] = 8'h10 ;
            rom[181] = 8'hd8 ;
            rom[182] = 8'hd1 ;
            rom[183] = 8'hf0 ;
            rom[184] = 8'h0c ;
            rom[185] = 8'h05 ;
            rom[186] = 8'hcc ;
            rom[187] = 8'he9 ;
            rom[188] = 8'h04 ;
            rom[189] = 8'h00 ;
            rom[190] = 8'hc6 ;
            rom[191] = 8'h0f ;
            rom[192] = 8'hed ;
            rom[193] = 8'hee ;
            rom[194] = 8'he0 ;
            rom[195] = 8'h09 ;
            rom[196] = 8'hfa ;
            rom[197] = 8'hfd ;
            rom[198] = 8'hf7 ;
            rom[199] = 8'hfe ;
            rom[200] = 8'hee ;
            rom[201] = 8'h30 ;
            rom[202] = 8'h05 ;
            rom[203] = 8'h00 ;
            rom[204] = 8'he4 ;
            rom[205] = 8'hf3 ;
            rom[206] = 8'h16 ;
            rom[207] = 8'hfb ;
            rom[208] = 8'hf9 ;
            rom[209] = 8'h11 ;
            rom[210] = 8'hbb ;
            rom[211] = 8'h02 ;
            rom[212] = 8'he5 ;
            rom[213] = 8'hea ;
            rom[214] = 8'h05 ;
            rom[215] = 8'h08 ;
            rom[216] = 8'hda ;
            rom[217] = 8'he9 ;
            rom[218] = 8'hc8 ;
            rom[219] = 8'he9 ;
            rom[220] = 8'he0 ;
            rom[221] = 8'h0e ;
            rom[222] = 8'h11 ;
            rom[223] = 8'h07 ;
            rom[224] = 8'he5 ;
            rom[225] = 8'hde ;
            rom[226] = 8'hf5 ;
            rom[227] = 8'hfc ;
            rom[228] = 8'hee ;
            rom[229] = 8'h13 ;
            rom[230] = 8'hde ;
            rom[231] = 8'hf3 ;
            rom[232] = 8'h01 ;
            rom[233] = 8'hf7 ;
            rom[234] = 8'he3 ;
            rom[235] = 8'he3 ;
            rom[236] = 8'h07 ;
            rom[237] = 8'hfc ;
            rom[238] = 8'hf7 ;
            rom[239] = 8'h01 ;
            rom[240] = 8'hcf ;
            rom[241] = 8'hc3 ;
            rom[242] = 8'he0 ;
            rom[243] = 8'h00 ;
            rom[244] = 8'hdc ;
            rom[245] = 8'h09 ;
            rom[246] = 8'hf2 ;
            rom[247] = 8'hdd ;
            rom[248] = 8'hf2 ;
            rom[249] = 8'h0d ;
            rom[250] = 8'h04 ;
            rom[251] = 8'h07 ;
            rom[252] = 8'h15 ;
            rom[253] = 8'hd0 ;
            rom[254] = 8'hb7 ;
            rom[255] = 8'he6 ;
            rom[256] = 8'h02 ;
            rom[257] = 8'hf8 ;
            rom[258] = 8'hd6 ;
            rom[259] = 8'h0e ;
            rom[260] = 8'h0e ;
            rom[261] = 8'hec ;
            rom[262] = 8'hff ;
            rom[263] = 8'hd2 ;
            rom[264] = 8'h06 ;
            rom[265] = 8'h1a ;
            rom[266] = 8'he0 ;
            rom[267] = 8'hec ;
            rom[268] = 8'he4 ;
            rom[269] = 8'h16 ;
            rom[270] = 8'h09 ;
            rom[271] = 8'h0b ;
            rom[272] = 8'h0d ;
            rom[273] = 8'h2f ;
            rom[274] = 8'hd4 ;
            rom[275] = 8'heb ;
            rom[276] = 8'h24 ;
            rom[277] = 8'h0b ;
            rom[278] = 8'hf6 ;
            rom[279] = 8'h1c ;
            rom[280] = 8'h1a ;
            rom[281] = 8'h17 ;
            rom[282] = 8'h06 ;
            rom[283] = 8'hff ;
            rom[284] = 8'h05 ;
            rom[285] = 8'h2a ;
            rom[286] = 8'h04 ;
            rom[287] = 8'h14 ;
            rom[288] = 8'hfa ;
            rom[289] = 8'h02 ;
            rom[290] = 8'hef ;
            rom[291] = 8'he6 ;
            rom[292] = 8'hf2 ;
            rom[293] = 8'h91 ;
            rom[294] = 8'he9 ;
            rom[295] = 8'h0a ;
            rom[296] = 8'he5 ;
            rom[297] = 8'hfa ;
            rom[298] = 8'hdf ;
            rom[299] = 8'hf3 ;
            rom[300] = 8'he5 ;
            rom[301] = 8'hc3 ;
            rom[302] = 8'h05 ;
            rom[303] = 8'he2 ;
            rom[304] = 8'he8 ;
            rom[305] = 8'hfd ;
            rom[306] = 8'hf3 ;
            rom[307] = 8'hfb ;
            rom[308] = 8'hff ;
            rom[309] = 8'hf3 ;
            rom[310] = 8'hc3 ;
            rom[311] = 8'hf2 ;
            rom[312] = 8'h38 ;
            rom[313] = 8'he2 ;
            rom[314] = 8'h00 ;
            rom[315] = 8'h04 ;
            rom[316] = 8'h0c ;
            rom[317] = 8'haa ;
            rom[318] = 8'h0b ;
            rom[319] = 8'he3 ;
            rom[320] = 8'hfd ;
            rom[321] = 8'h0d ;
            rom[322] = 8'hf1 ;
            rom[323] = 8'h05 ;
            rom[324] = 8'h11 ;
            rom[325] = 8'hab ;
            rom[326] = 8'h02 ;
            rom[327] = 8'h08 ;
            rom[328] = 8'hf3 ;
            rom[329] = 8'hfd ;
            rom[330] = 8'h0c ;
            rom[331] = 8'h1d ;
            rom[332] = 8'h08 ;
            rom[333] = 8'h0a ;
            rom[334] = 8'he0 ;
            rom[335] = 8'h0d ;
            rom[336] = 8'he0 ;
            rom[337] = 8'hf4 ;
            rom[338] = 8'h17 ;
            rom[339] = 8'h13 ;
            rom[340] = 8'h02 ;
            rom[341] = 8'h22 ;
            rom[342] = 8'hfe ;
            rom[343] = 8'h03 ;
            rom[344] = 8'hf9 ;
            rom[345] = 8'h0a ;
            rom[346] = 8'hf3 ;
            rom[347] = 8'hf8 ;
            rom[348] = 8'h15 ;
            rom[349] = 8'h1d ;
            rom[350] = 8'hef ;
            rom[351] = 8'hf5 ;
            rom[352] = 8'h0a ;
            rom[353] = 8'h03 ;
            rom[354] = 8'h12 ;
            rom[355] = 8'hbc ;
            rom[356] = 8'hcb ;
            rom[357] = 8'hd5 ;
            rom[358] = 8'hf0 ;
            rom[359] = 8'hfa ;
            rom[360] = 8'hf0 ;
            rom[361] = 8'hef ;
            rom[362] = 8'hda ;
            rom[363] = 8'hf3 ;
            rom[364] = 8'h05 ;
            rom[365] = 8'hc9 ;
            rom[366] = 8'hf9 ;
            rom[367] = 8'h17 ;
            rom[368] = 8'hff ;
            rom[369] = 8'h05 ;
            rom[370] = 8'hf6 ;
            rom[371] = 8'h15 ;
            rom[372] = 8'h0a ;
            rom[373] = 8'hd9 ;
            rom[374] = 8'h06 ;
            rom[375] = 8'hfe ;
            rom[376] = 8'hf1 ;
            rom[377] = 8'h14 ;
            rom[378] = 8'hf1 ;
            rom[379] = 8'hf8 ;
            rom[380] = 8'h09 ;
            rom[381] = 8'hec ;
            rom[382] = 8'hda ;
            rom[383] = 8'hff ;
            rom[384] = 8'hc3 ;
            rom[385] = 8'h00 ;
            rom[386] = 8'h26 ;
            rom[387] = 8'h1e ;
            rom[388] = 8'he4 ;
            rom[389] = 8'hf2 ;
            rom[390] = 8'h30 ;
            rom[391] = 8'h13 ;
            rom[392] = 8'hdf ;
            rom[393] = 8'hf8 ;
            rom[394] = 8'hcf ;
            rom[395] = 8'hde ;
            rom[396] = 8'hd3 ;
            rom[397] = 8'hf7 ;
            rom[398] = 8'hf1 ;
            rom[399] = 8'h0f ;
            rom[400] = 8'h11 ;
            rom[401] = 8'hfc ;
            rom[402] = 8'hd9 ;
            rom[403] = 8'hee ;
            rom[404] = 8'h12 ;
            rom[405] = 8'hdc ;
            rom[406] = 8'h02 ;
            rom[407] = 8'hf7 ;
            rom[408] = 8'hfd ;
            rom[409] = 8'hf0 ;
            rom[410] = 8'h07 ;
            rom[411] = 8'hf4 ;
            rom[412] = 8'h0d ;
            rom[413] = 8'hf8 ;
            rom[414] = 8'hf2 ;
            rom[415] = 8'hc7 ;
            rom[416] = 8'hfa ;
            rom[417] = 8'hfe ;
            rom[418] = 8'h2a ;
            rom[419] = 8'hfc ;
            rom[420] = 8'hff ;
            rom[421] = 8'h0a ;
            rom[422] = 8'hea ;
            rom[423] = 8'he3 ;
            rom[424] = 8'hec ;
            rom[425] = 8'he3 ;
            rom[426] = 8'h0b ;
            rom[427] = 8'hfe ;
            rom[428] = 8'h05 ;
            rom[429] = 8'h10 ;
            rom[430] = 8'h02 ;
            rom[431] = 8'hf0 ;
            rom[432] = 8'h1d ;
            rom[433] = 8'h12 ;
            rom[434] = 8'hf9 ;
            rom[435] = 8'h1f ;
            rom[436] = 8'hf7 ;
            rom[437] = 8'hf9 ;
            rom[438] = 8'hd7 ;
            rom[439] = 8'hda ;
            rom[440] = 8'hf8 ;
            rom[441] = 8'hff ;
            rom[442] = 8'hf0 ;
            rom[443] = 8'h0e ;
            rom[444] = 8'hf1 ;
            rom[445] = 8'hf4 ;
            rom[446] = 8'he0 ;
            rom[447] = 8'h0a ;
            rom[448] = 8'h0b ;
            rom[449] = 8'hee ;
            rom[450] = 8'hdc ;
            rom[451] = 8'hce ;
            rom[452] = 8'hc9 ;
            rom[453] = 8'hbd ;
            rom[454] = 8'he4 ;
            rom[455] = 8'hf9 ;
            rom[456] = 8'hd4 ;
            rom[457] = 8'hf3 ;
            rom[458] = 8'h1a ;
            rom[459] = 8'h2d ;
            rom[460] = 8'h00 ;
            rom[461] = 8'h0d ;
            rom[462] = 8'he7 ;
            rom[463] = 8'h0b ;
            rom[464] = 8'hf9 ;
            rom[465] = 8'hf8 ;
            rom[466] = 8'hcd ;
            rom[467] = 8'hed ;
            rom[468] = 8'h0d ;
            rom[469] = 8'hfb ;
            rom[470] = 8'hef ;
            rom[471] = 8'hf1 ;
            rom[472] = 8'h2e ;
            rom[473] = 8'h10 ;
            rom[474] = 8'h0f ;
            rom[475] = 8'hda ;
            rom[476] = 8'hed ;
            rom[477] = 8'h15 ;
            rom[478] = 8'hd8 ;
            rom[479] = 8'hf8 ;
            rom[480] = 8'hf7 ;
            rom[481] = 8'h13 ;
            rom[482] = 8'h05 ;
            rom[483] = 8'hfb ;
            rom[484] = 8'h21 ;
            rom[485] = 8'hf7 ;
            rom[486] = 8'h03 ;
            rom[487] = 8'hfc ;
            rom[488] = 8'hec ;
            rom[489] = 8'hed ;
            rom[490] = 8'hfe ;
            rom[491] = 8'hdb ;
            rom[492] = 8'hde ;
            rom[493] = 8'he0 ;
            rom[494] = 8'hff ;
            rom[495] = 8'h06 ;
            rom[496] = 8'h01 ;
            rom[497] = 8'h00 ;
            rom[498] = 8'h19 ;
            rom[499] = 8'hc1 ;
            rom[500] = 8'h06 ;
            rom[501] = 8'he5 ;
            rom[502] = 8'h09 ;
            rom[503] = 8'h0e ;
            rom[504] = 8'hf6 ;
            rom[505] = 8'hf2 ;
            rom[506] = 8'h1d ;
            rom[507] = 8'he4 ;
            rom[508] = 8'hed ;
            rom[509] = 8'hb0 ;
            rom[510] = 8'hef ;
            rom[511] = 8'hfc ;
            rom[512] = 8'h08 ;
            rom[513] = 8'hfe ;
            rom[514] = 8'hf5 ;
            rom[515] = 8'h1e ;
            rom[516] = 8'h03 ;
            rom[517] = 8'h07 ;
            rom[518] = 8'h05 ;
            rom[519] = 8'hfd ;
            rom[520] = 8'hf8 ;
            rom[521] = 8'hfa ;
            rom[522] = 8'hf8 ;
            rom[523] = 8'hdf ;
            rom[524] = 8'hef ;
            rom[525] = 8'h0b ;
            rom[526] = 8'h04 ;
            rom[527] = 8'hce ;
            rom[528] = 8'hb5 ;
            rom[529] = 8'hfe ;
            rom[530] = 8'hea ;
            rom[531] = 8'hf5 ;
            rom[532] = 8'hd6 ;
            rom[533] = 8'h02 ;
            rom[534] = 8'h03 ;
            rom[535] = 8'h09 ;
            rom[536] = 8'hff ;
            rom[537] = 8'hfb ;
            rom[538] = 8'he9 ;
            rom[539] = 8'h04 ;
            rom[540] = 8'h15 ;
            rom[541] = 8'h00 ;
            rom[542] = 8'h04 ;
            rom[543] = 8'h0b ;
            rom[544] = 8'h12 ;
            rom[545] = 8'h03 ;
            rom[546] = 8'h01 ;
            rom[547] = 8'hf8 ;
            rom[548] = 8'hde ;
            rom[549] = 8'he9 ;
            rom[550] = 8'h1b ;
            rom[551] = 8'h24 ;
            rom[552] = 8'hf5 ;
            rom[553] = 8'hfa ;
            rom[554] = 8'h10 ;
            rom[555] = 8'h18 ;
            rom[556] = 8'heb ;
            rom[557] = 8'he0 ;
            rom[558] = 8'hde ;
            rom[559] = 8'h14 ;
            rom[560] = 8'hd4 ;
            rom[561] = 8'hfc ;
            rom[562] = 8'hf0 ;
            rom[563] = 8'he5 ;
            rom[564] = 8'hee ;
            rom[565] = 8'h08 ;
            rom[566] = 8'he2 ;
            rom[567] = 8'h09 ;
            rom[568] = 8'h0f ;
            rom[569] = 8'h08 ;
            rom[570] = 8'h03 ;
            rom[571] = 8'hf0 ;
            rom[572] = 8'h0c ;
            rom[573] = 8'h0d ;
            rom[574] = 8'hef ;
            rom[575] = 8'he8 ;
            rom[576] = 8'hf3 ;
            rom[577] = 8'hfa ;
            rom[578] = 8'h18 ;
            rom[579] = 8'hfe ;
            rom[580] = 8'h19 ;
            rom[581] = 8'h0d ;
            rom[582] = 8'he7 ;
            rom[583] = 8'hd6 ;
            rom[584] = 8'hf8 ;
            rom[585] = 8'hfe ;
            rom[586] = 8'he3 ;
            rom[587] = 8'hed ;
            rom[588] = 8'hdd ;
            rom[589] = 8'h0e ;
            rom[590] = 8'hd8 ;
            rom[591] = 8'hf4 ;
            rom[592] = 8'hde ;
            rom[593] = 8'h16 ;
            rom[594] = 8'h04 ;
            rom[595] = 8'h07 ;
            rom[596] = 8'hfa ;
            rom[597] = 8'hf7 ;
            rom[598] = 8'hf6 ;
            rom[599] = 8'hda ;
            rom[600] = 8'hd4 ;
            rom[601] = 8'hf5 ;
            rom[602] = 8'hda ;
            rom[603] = 8'he2 ;
            rom[604] = 8'h08 ;
            rom[605] = 8'h1c ;
            rom[606] = 8'h25 ;
            rom[607] = 8'he3 ;
            rom[608] = 8'hff ;
            rom[609] = 8'hf5 ;
            rom[610] = 8'he1 ;
            rom[611] = 8'h12 ;
            rom[612] = 8'hc9 ;
            rom[613] = 8'h0b ;
            rom[614] = 8'hf5 ;
            rom[615] = 8'he2 ;
            rom[616] = 8'hed ;
            rom[617] = 8'h12 ;
            rom[618] = 8'h20 ;
            rom[619] = 8'h0a ;
            rom[620] = 8'hde ;
            rom[621] = 8'he1 ;
            rom[622] = 8'hfc ;
            rom[623] = 8'h00 ;
            rom[624] = 8'heb ;
            rom[625] = 8'h09 ;
            rom[626] = 8'h1e ;
            rom[627] = 8'h03 ;
            rom[628] = 8'hf0 ;
            rom[629] = 8'h0c ;
            rom[630] = 8'hf8 ;
            rom[631] = 8'h01 ;
            rom[632] = 8'he3 ;
            rom[633] = 8'hfa ;
            rom[634] = 8'hd9 ;
            rom[635] = 8'h04 ;
            rom[636] = 8'he0 ;
            rom[637] = 8'h29 ;
            rom[638] = 8'h08 ;
            rom[639] = 8'hdd ;
            rom[640] = 8'h01 ;
            rom[641] = 8'h0a ;
            rom[642] = 8'h0a ;
            rom[643] = 8'h11 ;
            rom[644] = 8'h10 ;
            rom[645] = 8'hdf ;
            rom[646] = 8'hf7 ;
            rom[647] = 8'h10 ;
            rom[648] = 8'he7 ;
            rom[649] = 8'h05 ;
            rom[650] = 8'h06 ;
            rom[651] = 8'h15 ;
            rom[652] = 8'hf2 ;
            rom[653] = 8'h19 ;
            rom[654] = 8'hd9 ;
            rom[655] = 8'h09 ;
            rom[656] = 8'h15 ;
            rom[657] = 8'hdb ;
            rom[658] = 8'h06 ;
            rom[659] = 8'hf1 ;
            rom[660] = 8'h03 ;
            rom[661] = 8'h0c ;
            rom[662] = 8'h05 ;
            rom[663] = 8'h16 ;
            rom[664] = 8'h23 ;
            rom[665] = 8'hfd ;
            rom[666] = 8'h1b ;
            rom[667] = 8'h21 ;
            rom[668] = 8'he2 ;
            rom[669] = 8'h1e ;
            rom[670] = 8'h0e ;
            rom[671] = 8'h25 ;
            rom[672] = 8'h05 ;
            rom[673] = 8'h07 ;
            rom[674] = 8'hef ;
            rom[675] = 8'h19 ;
            rom[676] = 8'hed ;
            rom[677] = 8'h29 ;
            rom[678] = 8'hd7 ;
            rom[679] = 8'h23 ;
            rom[680] = 8'h0a ;
            rom[681] = 8'h18 ;
            rom[682] = 8'h13 ;
            rom[683] = 8'hda ;
            rom[684] = 8'he4 ;
            rom[685] = 8'h1d ;
            rom[686] = 8'hfe ;
            rom[687] = 8'hfe ;
            rom[688] = 8'h05 ;
            rom[689] = 8'h18 ;
            rom[690] = 8'he0 ;
            rom[691] = 8'hf7 ;
            rom[692] = 8'h0a ;
            rom[693] = 8'hd6 ;
            rom[694] = 8'h09 ;
            rom[695] = 8'h4e ;
            rom[696] = 8'h26 ;
            rom[697] = 8'hf2 ;
            rom[698] = 8'h1b ;
            rom[699] = 8'hd6 ;
            rom[700] = 8'hf4 ;
            rom[701] = 8'hd3 ;
            rom[702] = 8'he7 ;
            rom[703] = 8'hf3 ;
            rom[704] = 8'hee ;
            rom[705] = 8'h04 ;
            rom[706] = 8'h13 ;
            rom[707] = 8'hf9 ;
            rom[708] = 8'h04 ;
            rom[709] = 8'he9 ;
            rom[710] = 8'heb ;
            rom[711] = 8'he5 ;
            rom[712] = 8'h00 ;
            rom[713] = 8'hf0 ;
            rom[714] = 8'h1f ;
            rom[715] = 8'h0f ;
            rom[716] = 8'h0e ;
            rom[717] = 8'h10 ;
            rom[718] = 8'hf3 ;
            rom[719] = 8'he8 ;
            rom[720] = 8'hf9 ;
            rom[721] = 8'h04 ;
            rom[722] = 8'h1d ;
            rom[723] = 8'h0a ;
            rom[724] = 8'hf8 ;
            rom[725] = 8'h0e ;
            rom[726] = 8'he6 ;
            rom[727] = 8'h03 ;
            rom[728] = 8'hee ;
            rom[729] = 8'h21 ;
            rom[730] = 8'h03 ;
            rom[731] = 8'hf2 ;
            rom[732] = 8'h0b ;
            rom[733] = 8'hf0 ;
            rom[734] = 8'hd2 ;
            rom[735] = 8'h09 ;
            rom[736] = 8'h08 ;
            rom[737] = 8'hfa ;
            rom[738] = 8'h17 ;
            rom[739] = 8'h02 ;
            rom[740] = 8'h07 ;
            rom[741] = 8'hee ;
            rom[742] = 8'hed ;
            rom[743] = 8'hf8 ;
            rom[744] = 8'he7 ;
            rom[745] = 8'hfc ;
            rom[746] = 8'hfa ;
            rom[747] = 8'hdc ;
            rom[748] = 8'he7 ;
            rom[749] = 8'h08 ;
            rom[750] = 8'h22 ;
            rom[751] = 8'h0e ;
            rom[752] = 8'h08 ;
            rom[753] = 8'h12 ;
            rom[754] = 8'h03 ;
            rom[755] = 8'h24 ;
            rom[756] = 8'he9 ;
            rom[757] = 8'h22 ;
            rom[758] = 8'h03 ;
            rom[759] = 8'hcf ;
            rom[760] = 8'hf3 ;
            rom[761] = 8'h13 ;
            rom[762] = 8'hfd ;
            rom[763] = 8'h0e ;
            rom[764] = 8'hf3 ;
            rom[765] = 8'heb ;
            rom[766] = 8'h10 ;
            rom[767] = 8'h1e ;
            rom[768] = 8'h02 ;
            rom[769] = 8'hc6 ;
            rom[770] = 8'h0b ;
            rom[771] = 8'hd8 ;
            rom[772] = 8'hda ;
            rom[773] = 8'hfb ;
            rom[774] = 8'hf7 ;
            rom[775] = 8'hd8 ;
            rom[776] = 8'h05 ;
            rom[777] = 8'hb9 ;
            rom[778] = 8'he5 ;
            rom[779] = 8'h1f ;
            rom[780] = 8'he8 ;
            rom[781] = 8'hd3 ;
            rom[782] = 8'h0a ;
            rom[783] = 8'hd8 ;
            rom[784] = 8'h0e ;
            rom[785] = 8'h02 ;
            rom[786] = 8'hf8 ;
            rom[787] = 8'h14 ;
            rom[788] = 8'hd7 ;
            rom[789] = 8'he9 ;
            rom[790] = 8'hf7 ;
            rom[791] = 8'h1d ;
            rom[792] = 8'hfd ;
            rom[793] = 8'hd3 ;
            rom[794] = 8'h0a ;
            rom[795] = 8'hc5 ;
            rom[796] = 8'h06 ;
            rom[797] = 8'he2 ;
            rom[798] = 8'heb ;
            rom[799] = 8'h25 ;
            rom[800] = 8'hf0 ;
            rom[801] = 8'h1d ;
            rom[802] = 8'h00 ;
            rom[803] = 8'hfc ;
            rom[804] = 8'h18 ;
            rom[805] = 8'h09 ;
            rom[806] = 8'h02 ;
            rom[807] = 8'hcf ;
            rom[808] = 8'h02 ;
            rom[809] = 8'heb ;
            rom[810] = 8'h11 ;
            rom[811] = 8'hfb ;
            rom[812] = 8'he2 ;
            rom[813] = 8'hf9 ;
            rom[814] = 8'h15 ;
            rom[815] = 8'hfb ;
            rom[816] = 8'hd1 ;
            rom[817] = 8'hfc ;
            rom[818] = 8'hdd ;
            rom[819] = 8'hfe ;
            rom[820] = 8'h0d ;
            rom[821] = 8'hef ;
            rom[822] = 8'hf3 ;
            rom[823] = 8'h10 ;
            rom[824] = 8'hfb ;
            rom[825] = 8'hf6 ;
            rom[826] = 8'hc6 ;
            rom[827] = 8'h0f ;
            rom[828] = 8'h25 ;
            rom[829] = 8'h09 ;
            rom[830] = 8'h0d ;
            rom[831] = 8'hc0 ;
            rom[832] = 8'hd5 ;
            rom[833] = 8'hfb ;
            rom[834] = 8'hfd ;
            rom[835] = 8'h17 ;
            rom[836] = 8'hfb ;
            rom[837] = 8'h29 ;
            rom[838] = 8'h10 ;
            rom[839] = 8'he7 ;
            rom[840] = 8'hf4 ;
            rom[841] = 8'hf6 ;
            rom[842] = 8'hea ;
            rom[843] = 8'hf9 ;
            rom[844] = 8'hd3 ;
            rom[845] = 8'hf4 ;
            rom[846] = 8'h12 ;
            rom[847] = 8'h12 ;
            rom[848] = 8'hd8 ;
            rom[849] = 8'h00 ;
            rom[850] = 8'h1d ;
            rom[851] = 8'hbe ;
            rom[852] = 8'heb ;
            rom[853] = 8'h10 ;
            rom[854] = 8'hee ;
            rom[855] = 8'h35 ;
            rom[856] = 8'hf3 ;
            rom[857] = 8'h1e ;
            rom[858] = 8'hef ;
            rom[859] = 8'h02 ;
            rom[860] = 8'hd9 ;
            rom[861] = 8'he1 ;
            rom[862] = 8'h13 ;
            rom[863] = 8'hef ;
            rom[864] = 8'h03 ;
            rom[865] = 8'hff ;
            rom[866] = 8'hcd ;
            rom[867] = 8'h13 ;
            rom[868] = 8'hd1 ;
            rom[869] = 8'h0c ;
            rom[870] = 8'h07 ;
            rom[871] = 8'h06 ;
            rom[872] = 8'he9 ;
            rom[873] = 8'hf5 ;
            rom[874] = 8'h09 ;
            rom[875] = 8'hfd ;
            rom[876] = 8'h20 ;
            rom[877] = 8'h14 ;
            rom[878] = 8'he1 ;
            rom[879] = 8'hef ;
            rom[880] = 8'hf2 ;
            rom[881] = 8'h04 ;
            rom[882] = 8'h1e ;
            rom[883] = 8'h0c ;
            rom[884] = 8'hf5 ;
            rom[885] = 8'h11 ;
            rom[886] = 8'h0e ;
            rom[887] = 8'he4 ;
            rom[888] = 8'h17 ;
            rom[889] = 8'hf2 ;
            rom[890] = 8'hd8 ;
            rom[891] = 8'h04 ;
            rom[892] = 8'h1c ;
            rom[893] = 8'hfb ;
            rom[894] = 8'hfe ;
            rom[895] = 8'h00 ;
            rom[896] = 8'h0f ;
            rom[897] = 8'hcb ;
            rom[898] = 8'heb ;
            rom[899] = 8'h32 ;
            rom[900] = 8'hf1 ;
            rom[901] = 8'he7 ;
            rom[902] = 8'h04 ;
            rom[903] = 8'hff ;
            rom[904] = 8'hde ;
            rom[905] = 8'hf2 ;
            rom[906] = 8'h05 ;
            rom[907] = 8'he6 ;
            rom[908] = 8'h01 ;
            rom[909] = 8'he9 ;
            rom[910] = 8'h05 ;
            rom[911] = 8'hf3 ;
            rom[912] = 8'h05 ;
            rom[913] = 8'hcd ;
            rom[914] = 8'he9 ;
            rom[915] = 8'h09 ;
            rom[916] = 8'h22 ;
            rom[917] = 8'hd7 ;
            rom[918] = 8'hd6 ;
            rom[919] = 8'hf9 ;
            rom[920] = 8'hce ;
            rom[921] = 8'h05 ;
            rom[922] = 8'hf3 ;
            rom[923] = 8'hd9 ;
            rom[924] = 8'h3a ;
            rom[925] = 8'h20 ;
            rom[926] = 8'h0e ;
            rom[927] = 8'h09 ;
            rom[928] = 8'h0f ;
            rom[929] = 8'h0a ;
            rom[930] = 8'hdd ;
            rom[931] = 8'hde ;
            rom[932] = 8'hdf ;
            rom[933] = 8'he8 ;
            rom[934] = 8'h05 ;
            rom[935] = 8'h02 ;
            rom[936] = 8'h01 ;
            rom[937] = 8'h17 ;
            rom[938] = 8'h36 ;
            rom[939] = 8'he9 ;
            rom[940] = 8'h1d ;
            rom[941] = 8'hf8 ;
            rom[942] = 8'he8 ;
            rom[943] = 8'h38 ;
            rom[944] = 8'h11 ;
            rom[945] = 8'h13 ;
            rom[946] = 8'hdf ;
            rom[947] = 8'hf5 ;
            rom[948] = 8'h11 ;
            rom[949] = 8'hfc ;
            rom[950] = 8'hf3 ;
            rom[951] = 8'h13 ;
            rom[952] = 8'hd1 ;
            rom[953] = 8'h15 ;
            rom[954] = 8'hf4 ;
            rom[955] = 8'hf9 ;
            rom[956] = 8'h22 ;
            rom[957] = 8'hf5 ;
            rom[958] = 8'hde ;
            rom[959] = 8'he4 ;
            rom[960] = 8'hfd ;
            rom[961] = 8'h27 ;
            rom[962] = 8'h03 ;
            rom[963] = 8'hf1 ;
            rom[964] = 8'h0a ;
            rom[965] = 8'hd5 ;
            rom[966] = 8'hf9 ;
            rom[967] = 8'h1a ;
            rom[968] = 8'h00 ;
            rom[969] = 8'h0d ;
            rom[970] = 8'hed ;
            rom[971] = 8'hf6 ;
            rom[972] = 8'hff ;
            rom[973] = 8'hf6 ;
            rom[974] = 8'hf4 ;
            rom[975] = 8'h29 ;
            rom[976] = 8'h1a ;
            rom[977] = 8'hf9 ;
            rom[978] = 8'he1 ;
            rom[979] = 8'h0c ;
            rom[980] = 8'hf9 ;
            rom[981] = 8'he2 ;
            rom[982] = 8'h20 ;
            rom[983] = 8'h40 ;
            rom[984] = 8'hf5 ;
            rom[985] = 8'h1e ;
            rom[986] = 8'h17 ;
            rom[987] = 8'hf7 ;
            rom[988] = 8'h8f ;
            rom[989] = 8'hcd ;
            rom[990] = 8'hfa ;
            rom[991] = 8'h05 ;
            rom[992] = 8'hf3 ;
            rom[993] = 8'h3b ;
            rom[994] = 8'hbe ;
            rom[995] = 8'he9 ;
            rom[996] = 8'he2 ;
            rom[997] = 8'h02 ;
            rom[998] = 8'h0a ;
            rom[999] = 8'he0 ;
            rom[1000] = 8'h0d ;
            rom[1001] = 8'h06 ;
            rom[1002] = 8'h0e ;
            rom[1003] = 8'hef ;
            rom[1004] = 8'h0e ;
            rom[1005] = 8'h09 ;
            rom[1006] = 8'hed ;
            rom[1007] = 8'hd8 ;
            rom[1008] = 8'h01 ;
            rom[1009] = 8'hfb ;
            rom[1010] = 8'hfd ;
            rom[1011] = 8'h16 ;
            rom[1012] = 8'h0e ;
            rom[1013] = 8'h14 ;
            rom[1014] = 8'he8 ;
            rom[1015] = 8'hf0 ;
            rom[1016] = 8'h01 ;
            rom[1017] = 8'hf5 ;
            rom[1018] = 8'he0 ;
            rom[1019] = 8'h07 ;
            rom[1020] = 8'hf0 ;
            rom[1021] = 8'h01 ;
            rom[1022] = 8'h1d ;
            rom[1023] = 8'hd7 ;
            rom[1024] = 8'hff ;
            rom[1025] = 8'h0f ;
            rom[1026] = 8'h1b ;
            rom[1027] = 8'h0f ;
            rom[1028] = 8'h04 ;
            rom[1029] = 8'hd6 ;
            rom[1030] = 8'h14 ;
            rom[1031] = 8'hf2 ;
            rom[1032] = 8'h03 ;
            rom[1033] = 8'h18 ;
            rom[1034] = 8'h09 ;
            rom[1035] = 8'h30 ;
            rom[1036] = 8'h09 ;
            rom[1037] = 8'heb ;
            rom[1038] = 8'hfe ;
            rom[1039] = 8'hdf ;
            rom[1040] = 8'hd0 ;
            rom[1041] = 8'h1f ;
            rom[1042] = 8'h00 ;
            rom[1043] = 8'hf3 ;
            rom[1044] = 8'h10 ;
            rom[1045] = 8'he5 ;
            rom[1046] = 8'hf4 ;
            rom[1047] = 8'hfd ;
            rom[1048] = 8'h04 ;
            rom[1049] = 8'hf9 ;
            rom[1050] = 8'h09 ;
            rom[1051] = 8'hd3 ;
            rom[1052] = 8'h23 ;
            rom[1053] = 8'h07 ;
            rom[1054] = 8'h08 ;
            rom[1055] = 8'h00 ;
            rom[1056] = 8'hf7 ;
            rom[1057] = 8'heb ;
            rom[1058] = 8'h07 ;
            rom[1059] = 8'h1e ;
            rom[1060] = 8'he4 ;
            rom[1061] = 8'hf3 ;
            rom[1062] = 8'h11 ;
            rom[1063] = 8'h0f ;
            rom[1064] = 8'hda ;
            rom[1065] = 8'hf8 ;
            rom[1066] = 8'heb ;
            rom[1067] = 8'hfc ;
            rom[1068] = 8'h05 ;
            rom[1069] = 8'hf3 ;
            rom[1070] = 8'heb ;
            rom[1071] = 8'hef ;
            rom[1072] = 8'hee ;
            rom[1073] = 8'h04 ;
            rom[1074] = 8'he4 ;
            rom[1075] = 8'hcc ;
            rom[1076] = 8'h25 ;
            rom[1077] = 8'hf1 ;
            rom[1078] = 8'hd0 ;
            rom[1079] = 8'hf0 ;
            rom[1080] = 8'h22 ;
            rom[1081] = 8'hea ;
            rom[1082] = 8'hf2 ;
            rom[1083] = 8'hf9 ;
            rom[1084] = 8'h03 ;
            rom[1085] = 8'h0d ;
            rom[1086] = 8'he4 ;
            rom[1087] = 8'hbe ;
            rom[1088] = 8'he0 ;
            rom[1089] = 8'h0e ;
            rom[1090] = 8'h26 ;
            rom[1091] = 8'h0d ;
            rom[1092] = 8'he1 ;
            rom[1093] = 8'hfe ;
            rom[1094] = 8'hd6 ;
            rom[1095] = 8'hef ;
            rom[1096] = 8'hf0 ;
            rom[1097] = 8'h15 ;
            rom[1098] = 8'hcd ;
            rom[1099] = 8'hda ;
            rom[1100] = 8'hf3 ;
            rom[1101] = 8'hd7 ;
            rom[1102] = 8'hea ;
            rom[1103] = 8'hfb ;
            rom[1104] = 8'h05 ;
            rom[1105] = 8'h19 ;
            rom[1106] = 8'hf6 ;
            rom[1107] = 8'h19 ;
            rom[1108] = 8'hfa ;
            rom[1109] = 8'he5 ;
            rom[1110] = 8'hea ;
            rom[1111] = 8'hd8 ;
            rom[1112] = 8'hd6 ;
            rom[1113] = 8'h04 ;
            rom[1114] = 8'he1 ;
            rom[1115] = 8'h27 ;
            rom[1116] = 8'h10 ;
            rom[1117] = 8'h0b ;
            rom[1118] = 8'h34 ;
            rom[1119] = 8'h08 ;
            rom[1120] = 8'hd2 ;
            rom[1121] = 8'hf8 ;
            rom[1122] = 8'hc9 ;
            rom[1123] = 8'h24 ;
            rom[1124] = 8'hf8 ;
            rom[1125] = 8'hf9 ;
            rom[1126] = 8'hcf ;
            rom[1127] = 8'he1 ;
            rom[1128] = 8'h16 ;
            rom[1129] = 8'h20 ;
            rom[1130] = 8'h07 ;
            rom[1131] = 8'hfe ;
            rom[1132] = 8'hf3 ;
            rom[1133] = 8'hf4 ;
            rom[1134] = 8'hd7 ;
            rom[1135] = 8'h0a ;
            rom[1136] = 8'hd6 ;
            rom[1137] = 8'hfa ;
            rom[1138] = 8'hfb ;
            rom[1139] = 8'hf7 ;
            rom[1140] = 8'hff ;
            rom[1141] = 8'hfe ;
            rom[1142] = 8'he8 ;
            rom[1143] = 8'heb ;
            rom[1144] = 8'hc4 ;
            rom[1145] = 8'hfa ;
            rom[1146] = 8'hee ;
            rom[1147] = 8'h0b ;
            rom[1148] = 8'hf6 ;
            rom[1149] = 8'h17 ;
            rom[1150] = 8'h14 ;
            rom[1151] = 8'he0 ;
            rom[1152] = 8'hf9 ;
            rom[1153] = 8'he2 ;
            rom[1154] = 8'h0e ;
            rom[1155] = 8'hed ;
            rom[1156] = 8'hf5 ;
            rom[1157] = 8'h03 ;
            rom[1158] = 8'h0d ;
            rom[1159] = 8'hc6 ;
            rom[1160] = 8'hf5 ;
            rom[1161] = 8'hea ;
            rom[1162] = 8'h04 ;
            rom[1163] = 8'h09 ;
            rom[1164] = 8'hf2 ;
            rom[1165] = 8'he1 ;
            rom[1166] = 8'h06 ;
            rom[1167] = 8'hd4 ;
            rom[1168] = 8'he4 ;
            rom[1169] = 8'hfd ;
            rom[1170] = 8'h1b ;
            rom[1171] = 8'h01 ;
            rom[1172] = 8'hf2 ;
            rom[1173] = 8'hee ;
            rom[1174] = 8'hec ;
            rom[1175] = 8'h09 ;
            rom[1176] = 8'hbf ;
            rom[1177] = 8'hec ;
            rom[1178] = 8'he4 ;
            rom[1179] = 8'hd8 ;
            rom[1180] = 8'hfb ;
            rom[1181] = 8'he4 ;
            rom[1182] = 8'hd1 ;
            rom[1183] = 8'h19 ;
            rom[1184] = 8'hee ;
            rom[1185] = 8'h11 ;
            rom[1186] = 8'h17 ;
            rom[1187] = 8'h1f ;
            rom[1188] = 8'h18 ;
            rom[1189] = 8'h01 ;
            rom[1190] = 8'h0c ;
            rom[1191] = 8'hce ;
            rom[1192] = 8'hfe ;
            rom[1193] = 8'h06 ;
            rom[1194] = 8'he9 ;
            rom[1195] = 8'h10 ;
            rom[1196] = 8'h33 ;
            rom[1197] = 8'h0a ;
            rom[1198] = 8'h19 ;
            rom[1199] = 8'hbf ;
            rom[1200] = 8'hec ;
            rom[1201] = 8'hba ;
            rom[1202] = 8'h0b ;
            rom[1203] = 8'hf4 ;
            rom[1204] = 8'h17 ;
            rom[1205] = 8'hc9 ;
            rom[1206] = 8'he0 ;
            rom[1207] = 8'h05 ;
            rom[1208] = 8'h10 ;
            rom[1209] = 8'h03 ;
            rom[1210] = 8'he8 ;
            rom[1211] = 8'hed ;
            rom[1212] = 8'h1c ;
            rom[1213] = 8'h05 ;
            rom[1214] = 8'h0c ;
            rom[1215] = 8'hf7 ;
            rom[1216] = 8'he5 ;
            rom[1217] = 8'hf4 ;
            rom[1218] = 8'h03 ;
            rom[1219] = 8'h0b ;
            rom[1220] = 8'he7 ;
            rom[1221] = 8'h01 ;
            rom[1222] = 8'h21 ;
            rom[1223] = 8'h06 ;
            rom[1224] = 8'heb ;
            rom[1225] = 8'h29 ;
            rom[1226] = 8'h0e ;
            rom[1227] = 8'hfa ;
            rom[1228] = 8'hdf ;
            rom[1229] = 8'h08 ;
            rom[1230] = 8'h0e ;
            rom[1231] = 8'h2e ;
            rom[1232] = 8'hd6 ;
            rom[1233] = 8'hef ;
            rom[1234] = 8'hfd ;
            rom[1235] = 8'h00 ;
            rom[1236] = 8'h0c ;
            rom[1237] = 8'h0f ;
            rom[1238] = 8'h14 ;
            rom[1239] = 8'hf5 ;
            rom[1240] = 8'hda ;
            rom[1241] = 8'hfe ;
            rom[1242] = 8'hd7 ;
            rom[1243] = 8'h11 ;
            rom[1244] = 8'hbe ;
            rom[1245] = 8'hf5 ;
            rom[1246] = 8'hfd ;
            rom[1247] = 8'h1e ;
            rom[1248] = 8'hf6 ;
            rom[1249] = 8'hdd ;
            rom[1250] = 8'h06 ;
            rom[1251] = 8'h02 ;
            rom[1252] = 8'hdb ;
            rom[1253] = 8'he0 ;
            rom[1254] = 8'hfb ;
            rom[1255] = 8'hf7 ;
            rom[1256] = 8'h06 ;
            rom[1257] = 8'hf3 ;
            rom[1258] = 8'h02 ;
            rom[1259] = 8'h0f ;
            rom[1260] = 8'h2b ;
            rom[1261] = 8'hd9 ;
            rom[1262] = 8'h12 ;
            rom[1263] = 8'hd8 ;
            rom[1264] = 8'hd4 ;
            rom[1265] = 8'hf6 ;
            rom[1266] = 8'h09 ;
            rom[1267] = 8'h16 ;
            rom[1268] = 8'h17 ;
            rom[1269] = 8'h04 ;
            rom[1270] = 8'hed ;
            rom[1271] = 8'h05 ;
            rom[1272] = 8'h11 ;
            rom[1273] = 8'he2 ;
            rom[1274] = 8'hfc ;
            rom[1275] = 8'h01 ;
            rom[1276] = 8'h1d ;
            rom[1277] = 8'hfc ;
            rom[1278] = 8'hf5 ;
            rom[1279] = 8'he6 ;
            rom[1280] = 8'hf8 ;
            rom[1281] = 8'hbf ;
            rom[1282] = 8'h00 ;
            rom[1283] = 8'h25 ;
            rom[1284] = 8'hdb ;
            rom[1285] = 8'hf9 ;
            rom[1286] = 8'h0f ;
            rom[1287] = 8'h00 ;
            rom[1288] = 8'hc7 ;
            rom[1289] = 8'h0a ;
            rom[1290] = 8'h1a ;
            rom[1291] = 8'hd9 ;
            rom[1292] = 8'h0b ;
            rom[1293] = 8'hd1 ;
            rom[1294] = 8'hfa ;
            rom[1295] = 8'hfa ;
            rom[1296] = 8'hd9 ;
            rom[1297] = 8'hcf ;
            rom[1298] = 8'hbb ;
            rom[1299] = 8'hf1 ;
            rom[1300] = 8'hf2 ;
            rom[1301] = 8'h00 ;
            rom[1302] = 8'h24 ;
            rom[1303] = 8'hf0 ;
            rom[1304] = 8'hfd ;
            rom[1305] = 8'he2 ;
            rom[1306] = 8'hf4 ;
            rom[1307] = 8'hf7 ;
            rom[1308] = 8'h06 ;
            rom[1309] = 8'h21 ;
            rom[1310] = 8'h09 ;
            rom[1311] = 8'h09 ;
            rom[1312] = 8'h0d ;
            rom[1313] = 8'he6 ;
            rom[1314] = 8'hd8 ;
            rom[1315] = 8'hf0 ;
            rom[1316] = 8'h21 ;
            rom[1317] = 8'hfe ;
            rom[1318] = 8'h02 ;
            rom[1319] = 8'h16 ;
            rom[1320] = 8'he2 ;
            rom[1321] = 8'h4c ;
            rom[1322] = 8'h0a ;
            rom[1323] = 8'he9 ;
            rom[1324] = 8'h1d ;
            rom[1325] = 8'h0d ;
            rom[1326] = 8'he5 ;
            rom[1327] = 8'hf0 ;
            rom[1328] = 8'h19 ;
            rom[1329] = 8'h20 ;
            rom[1330] = 8'h1f ;
            rom[1331] = 8'hfe ;
            rom[1332] = 8'hf6 ;
            rom[1333] = 8'h20 ;
            rom[1334] = 8'heb ;
            rom[1335] = 8'h08 ;
            rom[1336] = 8'h04 ;
            rom[1337] = 8'h04 ;
            rom[1338] = 8'hfd ;
            rom[1339] = 8'h04 ;
            rom[1340] = 8'h09 ;
            rom[1341] = 8'h11 ;
            rom[1342] = 8'he0 ;
            rom[1343] = 8'he6 ;
            rom[1344] = 8'h1a ;
            rom[1345] = 8'h06 ;
            rom[1346] = 8'h23 ;
            rom[1347] = 8'hc7 ;
            rom[1348] = 8'h07 ;
            rom[1349] = 8'hf3 ;
            rom[1350] = 8'hf5 ;
            rom[1351] = 8'hd7 ;
            rom[1352] = 8'h13 ;
            rom[1353] = 8'hfc ;
            rom[1354] = 8'hc7 ;
            rom[1355] = 8'h19 ;
            rom[1356] = 8'he9 ;
            rom[1357] = 8'h0b ;
            rom[1358] = 8'hec ;
            rom[1359] = 8'h1e ;
            rom[1360] = 8'h05 ;
            rom[1361] = 8'hf3 ;
            rom[1362] = 8'hed ;
            rom[1363] = 8'he0 ;
            rom[1364] = 8'h0e ;
            rom[1365] = 8'hef ;
            rom[1366] = 8'hf7 ;
            rom[1367] = 8'h0f ;
            rom[1368] = 8'hef ;
            rom[1369] = 8'h1d ;
            rom[1370] = 8'hf3 ;
            rom[1371] = 8'hed ;
            rom[1372] = 8'he6 ;
            rom[1373] = 8'he4 ;
            rom[1374] = 8'hc5 ;
            rom[1375] = 8'he9 ;
            rom[1376] = 8'hfc ;
            rom[1377] = 8'h17 ;
            rom[1378] = 8'h21 ;
            rom[1379] = 8'hfe ;
            rom[1380] = 8'hff ;
            rom[1381] = 8'heb ;
            rom[1382] = 8'h17 ;
            rom[1383] = 8'h01 ;
            rom[1384] = 8'hb6 ;
            rom[1385] = 8'h1a ;
            rom[1386] = 8'h0f ;
            rom[1387] = 8'hf8 ;
            rom[1388] = 8'he4 ;
            rom[1389] = 8'hdd ;
            rom[1390] = 8'h04 ;
            rom[1391] = 8'h09 ;
            rom[1392] = 8'h18 ;
            rom[1393] = 8'hf0 ;
            rom[1394] = 8'hea ;
            rom[1395] = 8'hf5 ;
            rom[1396] = 8'h0e ;
            rom[1397] = 8'he6 ;
            rom[1398] = 8'h0c ;
            rom[1399] = 8'heb ;
            rom[1400] = 8'h19 ;
            rom[1401] = 8'hf4 ;
            rom[1402] = 8'hfc ;
            rom[1403] = 8'h0f ;
            rom[1404] = 8'he9 ;
            rom[1405] = 8'hf7 ;
            rom[1406] = 8'heb ;
            rom[1407] = 8'h1c ;
            rom[1408] = 8'hff ;
            rom[1409] = 8'h03 ;
            rom[1410] = 8'hfd ;
            rom[1411] = 8'he4 ;
            rom[1412] = 8'he5 ;
            rom[1413] = 8'he3 ;
            rom[1414] = 8'hfb ;
            rom[1415] = 8'h03 ;
            rom[1416] = 8'hef ;
            rom[1417] = 8'h03 ;
            rom[1418] = 8'h06 ;
            rom[1419] = 8'hc3 ;
            rom[1420] = 8'hf4 ;
            rom[1421] = 8'hdc ;
            rom[1422] = 8'h16 ;
            rom[1423] = 8'hba ;
            rom[1424] = 8'h0c ;
            rom[1425] = 8'he9 ;
            rom[1426] = 8'he1 ;
            rom[1427] = 8'h02 ;
            rom[1428] = 8'h15 ;
            rom[1429] = 8'he5 ;
            rom[1430] = 8'h1b ;
            rom[1431] = 8'h11 ;
            rom[1432] = 8'h05 ;
            rom[1433] = 8'h01 ;
            rom[1434] = 8'hc3 ;
            rom[1435] = 8'he0 ;
            rom[1436] = 8'h0b ;
            rom[1437] = 8'hf9 ;
            rom[1438] = 8'h13 ;
            rom[1439] = 8'h05 ;
            rom[1440] = 8'hf7 ;
            rom[1441] = 8'h05 ;
            rom[1442] = 8'h03 ;
            rom[1443] = 8'hfe ;
            rom[1444] = 8'hfd ;
            rom[1445] = 8'hfc ;
            rom[1446] = 8'hee ;
            rom[1447] = 8'hf7 ;
            rom[1448] = 8'hf4 ;
            rom[1449] = 8'hf2 ;
            rom[1450] = 8'hdf ;
            rom[1451] = 8'hfe ;
            rom[1452] = 8'h0d ;
            rom[1453] = 8'he1 ;
            rom[1454] = 8'hde ;
            rom[1455] = 8'hf6 ;
            rom[1456] = 8'h1f ;
            rom[1457] = 8'h15 ;
            rom[1458] = 8'hd0 ;
            rom[1459] = 8'h16 ;
            rom[1460] = 8'hfb ;
            rom[1461] = 8'h00 ;
            rom[1462] = 8'h12 ;
            rom[1463] = 8'hc7 ;
            rom[1464] = 8'hf1 ;
            rom[1465] = 8'h1b ;
            rom[1466] = 8'h11 ;
            rom[1467] = 8'he1 ;
            rom[1468] = 8'h0a ;
            rom[1469] = 8'hf2 ;
            rom[1470] = 8'h00 ;
            rom[1471] = 8'he7 ;
            rom[1472] = 8'hfc ;
            rom[1473] = 8'hf7 ;
            rom[1474] = 8'h0c ;
            rom[1475] = 8'hee ;
            rom[1476] = 8'hf0 ;
            rom[1477] = 8'h10 ;
            rom[1478] = 8'hed ;
            rom[1479] = 8'hf4 ;
            rom[1480] = 8'h09 ;
            rom[1481] = 8'hfd ;
            rom[1482] = 8'hda ;
            rom[1483] = 8'hf1 ;
            rom[1484] = 8'hf6 ;
            rom[1485] = 8'h24 ;
            rom[1486] = 8'hf0 ;
            rom[1487] = 8'h23 ;
            rom[1488] = 8'h09 ;
            rom[1489] = 8'hd8 ;
            rom[1490] = 8'h18 ;
            rom[1491] = 8'he4 ;
            rom[1492] = 8'hdf ;
            rom[1493] = 8'hf7 ;
            rom[1494] = 8'hc0 ;
            rom[1495] = 8'h16 ;
            rom[1496] = 8'h0b ;
            rom[1497] = 8'hd4 ;
            rom[1498] = 8'h0e ;
            rom[1499] = 8'h25 ;
            rom[1500] = 8'h0a ;
            rom[1501] = 8'h0f ;
            rom[1502] = 8'hff ;
            rom[1503] = 8'hf4 ;
            rom[1504] = 8'h05 ;
            rom[1505] = 8'hfe ;
            rom[1506] = 8'heb ;
            rom[1507] = 8'h0d ;
            rom[1508] = 8'h05 ;
            rom[1509] = 8'hfd ;
            rom[1510] = 8'hea ;
            rom[1511] = 8'h05 ;
            rom[1512] = 8'hd0 ;
            rom[1513] = 8'hfd ;
            rom[1514] = 8'h0c ;
            rom[1515] = 8'h07 ;
            rom[1516] = 8'h20 ;
            rom[1517] = 8'h0c ;
            rom[1518] = 8'he9 ;
            rom[1519] = 8'hf3 ;
            rom[1520] = 8'h03 ;
            rom[1521] = 8'hd6 ;
            rom[1522] = 8'hff ;
            rom[1523] = 8'he9 ;
            rom[1524] = 8'hfe ;
            rom[1525] = 8'hf8 ;
            rom[1526] = 8'hce ;
            rom[1527] = 8'h0a ;
            rom[1528] = 8'hfe ;
            rom[1529] = 8'hbd ;
            rom[1530] = 8'hed ;
            rom[1531] = 8'h01 ;
            rom[1532] = 8'he6 ;
            rom[1533] = 8'h00 ;
            rom[1534] = 8'h0c ;
            rom[1535] = 8'hec ;
            rom[1536] = 8'hda ;
            rom[1537] = 8'hd9 ;
            rom[1538] = 8'h0d ;
            rom[1539] = 8'hcf ;
            rom[1540] = 8'h04 ;
            rom[1541] = 8'h16 ;
            rom[1542] = 8'hfb ;
            rom[1543] = 8'hf5 ;
            rom[1544] = 8'h00 ;
            rom[1545] = 8'he4 ;
            rom[1546] = 8'h0d ;
            rom[1547] = 8'he6 ;
            rom[1548] = 8'h29 ;
            rom[1549] = 8'hde ;
            rom[1550] = 8'h31 ;
            rom[1551] = 8'heb ;
            rom[1552] = 8'h1d ;
            rom[1553] = 8'ha9 ;
            rom[1554] = 8'h0a ;
            rom[1555] = 8'h33 ;
            rom[1556] = 8'hef ;
            rom[1557] = 8'he1 ;
            rom[1558] = 8'h15 ;
            rom[1559] = 8'h02 ;
            rom[1560] = 8'h32 ;
            rom[1561] = 8'he1 ;
            rom[1562] = 8'hfb ;
            rom[1563] = 8'h09 ;
            rom[1564] = 8'hed ;
            rom[1565] = 8'h0d ;
            rom[1566] = 8'h12 ;
            rom[1567] = 8'he7 ;
            rom[1568] = 8'hf1 ;
            rom[1569] = 8'hf2 ;
            rom[1570] = 8'h00 ;
            rom[1571] = 8'hcd ;
            rom[1572] = 8'h20 ;
            rom[1573] = 8'h15 ;
            rom[1574] = 8'hf7 ;
            rom[1575] = 8'hdc ;
            rom[1576] = 8'h2a ;
            rom[1577] = 8'hd5 ;
            rom[1578] = 8'h00 ;
            rom[1579] = 8'h1b ;
            rom[1580] = 8'hdd ;
            rom[1581] = 8'h27 ;
            rom[1582] = 8'he5 ;
            rom[1583] = 8'he2 ;
            rom[1584] = 8'h16 ;
            rom[1585] = 8'h14 ;
            rom[1586] = 8'h01 ;
            rom[1587] = 8'h03 ;
            rom[1588] = 8'heb ;
            rom[1589] = 8'h0f ;
            rom[1590] = 8'h21 ;
            rom[1591] = 8'hf9 ;
            rom[1592] = 8'hf2 ;
            rom[1593] = 8'h10 ;
            rom[1594] = 8'h02 ;
            rom[1595] = 8'hfe ;
            rom[1596] = 8'hfd ;
            rom[1597] = 8'h02 ;
            rom[1598] = 8'hef ;
            rom[1599] = 8'hfa ;
            rom[1600] = 8'h08 ;
            rom[1601] = 8'hcc ;
            rom[1602] = 8'hf4 ;
            rom[1603] = 8'h1b ;
            rom[1604] = 8'hdb ;
            rom[1605] = 8'h31 ;
            rom[1606] = 8'h00 ;
            rom[1607] = 8'he4 ;
            rom[1608] = 8'hdb ;
            rom[1609] = 8'hfd ;
            rom[1610] = 8'hc3 ;
            rom[1611] = 8'h05 ;
            rom[1612] = 8'hf7 ;
            rom[1613] = 8'h13 ;
            rom[1614] = 8'h16 ;
            rom[1615] = 8'he8 ;
            rom[1616] = 8'h12 ;
            rom[1617] = 8'he0 ;
            rom[1618] = 8'h0e ;
            rom[1619] = 8'hfb ;
            rom[1620] = 8'h2e ;
            rom[1621] = 8'h06 ;
            rom[1622] = 8'h07 ;
            rom[1623] = 8'hfb ;
            rom[1624] = 8'h08 ;
            rom[1625] = 8'hfe ;
            rom[1626] = 8'he6 ;
            rom[1627] = 8'hff ;
            rom[1628] = 8'h09 ;
            rom[1629] = 8'hf5 ;
            rom[1630] = 8'hde ;
            rom[1631] = 8'hd3 ;
            rom[1632] = 8'h1a ;
            rom[1633] = 8'h07 ;
            rom[1634] = 8'hd5 ;
            rom[1635] = 8'h00 ;
            rom[1636] = 8'h0f ;
            rom[1637] = 8'h31 ;
            rom[1638] = 8'hfc ;
            rom[1639] = 8'hee ;
            rom[1640] = 8'h08 ;
            rom[1641] = 8'hc9 ;
            rom[1642] = 8'hf5 ;
            rom[1643] = 8'h11 ;
            rom[1644] = 8'hf8 ;
            rom[1645] = 8'h12 ;
            rom[1646] = 8'hdd ;
            rom[1647] = 8'h03 ;
            rom[1648] = 8'hfe ;
            rom[1649] = 8'hf7 ;
            rom[1650] = 8'h25 ;
            rom[1651] = 8'hb3 ;
            rom[1652] = 8'h07 ;
            rom[1653] = 8'h1c ;
            rom[1654] = 8'he3 ;
            rom[1655] = 8'h01 ;
            rom[1656] = 8'h02 ;
            rom[1657] = 8'hd7 ;
            rom[1658] = 8'hff ;
            rom[1659] = 8'hf5 ;
            rom[1660] = 8'hec ;
            rom[1661] = 8'hf4 ;
            rom[1662] = 8'hee ;
            rom[1663] = 8'h1f ;
            rom[1664] = 8'he9 ;
            rom[1665] = 8'hfa ;
            rom[1666] = 8'he6 ;
            rom[1667] = 8'h0f ;
            rom[1668] = 8'h26 ;
            rom[1669] = 8'h11 ;
            rom[1670] = 8'hee ;
            rom[1671] = 8'h0b ;
            rom[1672] = 8'h0e ;
            rom[1673] = 8'hdd ;
            rom[1674] = 8'hfa ;
            rom[1675] = 8'h0c ;
            rom[1676] = 8'h09 ;
            rom[1677] = 8'hf8 ;
            rom[1678] = 8'h0f ;
            rom[1679] = 8'hf3 ;
            rom[1680] = 8'h01 ;
            rom[1681] = 8'h02 ;
            rom[1682] = 8'hf0 ;
            rom[1683] = 8'hff ;
            rom[1684] = 8'hf3 ;
            rom[1685] = 8'hf2 ;
            rom[1686] = 8'hfd ;
            rom[1687] = 8'h04 ;
            rom[1688] = 8'he1 ;
            rom[1689] = 8'hd1 ;
            rom[1690] = 8'h10 ;
            rom[1691] = 8'hee ;
            rom[1692] = 8'h0b ;
            rom[1693] = 8'he9 ;
            rom[1694] = 8'hf7 ;
            rom[1695] = 8'h01 ;
            rom[1696] = 8'h0e ;
            rom[1697] = 8'h29 ;
            rom[1698] = 8'hcf ;
            rom[1699] = 8'h0c ;
            rom[1700] = 8'hcf ;
            rom[1701] = 8'h11 ;
            rom[1702] = 8'he2 ;
            rom[1703] = 8'h19 ;
            rom[1704] = 8'h04 ;
            rom[1705] = 8'hea ;
            rom[1706] = 8'h0a ;
            rom[1707] = 8'h02 ;
            rom[1708] = 8'h09 ;
            rom[1709] = 8'hd3 ;
            rom[1710] = 8'hf6 ;
            rom[1711] = 8'hdf ;
            rom[1712] = 8'hed ;
            rom[1713] = 8'h27 ;
            rom[1714] = 8'hd4 ;
            rom[1715] = 8'hf4 ;
            rom[1716] = 8'hc8 ;
            rom[1717] = 8'h18 ;
            rom[1718] = 8'h1e ;
            rom[1719] = 8'h06 ;
            rom[1720] = 8'hff ;
            rom[1721] = 8'hc7 ;
            rom[1722] = 8'h26 ;
            rom[1723] = 8'hcd ;
            rom[1724] = 8'hec ;
            rom[1725] = 8'h09 ;
            rom[1726] = 8'hf8 ;
            rom[1727] = 8'hf3 ;
            rom[1728] = 8'h0f ;
            rom[1729] = 8'hf0 ;
            rom[1730] = 8'h06 ;
            rom[1731] = 8'he6 ;
            rom[1732] = 8'hff ;
            rom[1733] = 8'h06 ;
            rom[1734] = 8'h07 ;
            rom[1735] = 8'hf1 ;
            rom[1736] = 8'h42 ;
            rom[1737] = 8'hd4 ;
            rom[1738] = 8'hd9 ;
            rom[1739] = 8'he9 ;
            rom[1740] = 8'hf7 ;
            rom[1741] = 8'h04 ;
            rom[1742] = 8'he2 ;
            rom[1743] = 8'h29 ;
            rom[1744] = 8'h12 ;
            rom[1745] = 8'hf5 ;
            rom[1746] = 8'h12 ;
            rom[1747] = 8'h0e ;
            rom[1748] = 8'hf6 ;
            rom[1749] = 8'h04 ;
            rom[1750] = 8'h09 ;
            rom[1751] = 8'hf5 ;
            rom[1752] = 8'h08 ;
            rom[1753] = 8'h1a ;
            rom[1754] = 8'h1d ;
            rom[1755] = 8'h14 ;
            rom[1756] = 8'hf2 ;
            rom[1757] = 8'h09 ;
            rom[1758] = 8'hf4 ;
            rom[1759] = 8'h0b ;
            rom[1760] = 8'h0d ;
            rom[1761] = 8'h0f ;
            rom[1762] = 8'h11 ;
            rom[1763] = 8'hf8 ;
            rom[1764] = 8'hee ;
            rom[1765] = 8'he3 ;
            rom[1766] = 8'hfd ;
            rom[1767] = 8'hf2 ;
            rom[1768] = 8'h28 ;
            rom[1769] = 8'hfe ;
            rom[1770] = 8'hf8 ;
            rom[1771] = 8'hfa ;
            rom[1772] = 8'hfd ;
            rom[1773] = 8'hf3 ;
            rom[1774] = 8'h09 ;
            rom[1775] = 8'h01 ;
            rom[1776] = 8'hfc ;
            rom[1777] = 8'hd9 ;
            rom[1778] = 8'he8 ;
            rom[1779] = 8'hf1 ;
            rom[1780] = 8'he1 ;
            rom[1781] = 8'hf6 ;
            rom[1782] = 8'h11 ;
            rom[1783] = 8'hfd ;
            rom[1784] = 8'h17 ;
            rom[1785] = 8'h3c ;
            rom[1786] = 8'h0c ;
            rom[1787] = 8'h13 ;
            rom[1788] = 8'hda ;
            rom[1789] = 8'h03 ;
            rom[1790] = 8'h0f ;
            rom[1791] = 8'h06 ;
            rom[1792] = 8'h00 ;
            rom[1793] = 8'h0f ;
            rom[1794] = 8'hfe ;
            rom[1795] = 8'h1b ;
            rom[1796] = 8'h22 ;
            rom[1797] = 8'h04 ;
            rom[1798] = 8'hf7 ;
            rom[1799] = 8'hdf ;
            rom[1800] = 8'hf2 ;
            rom[1801] = 8'hff ;
            rom[1802] = 8'hf4 ;
            rom[1803] = 8'hd5 ;
            rom[1804] = 8'he4 ;
            rom[1805] = 8'h12 ;
            rom[1806] = 8'hfc ;
            rom[1807] = 8'h12 ;
            rom[1808] = 8'h11 ;
            rom[1809] = 8'h1b ;
            rom[1810] = 8'hda ;
            rom[1811] = 8'h0a ;
            rom[1812] = 8'hf5 ;
            rom[1813] = 8'hf1 ;
            rom[1814] = 8'hff ;
            rom[1815] = 8'h18 ;
            rom[1816] = 8'hff ;
            rom[1817] = 8'h08 ;
            rom[1818] = 8'h0c ;
            rom[1819] = 8'h09 ;
            rom[1820] = 8'hdd ;
            rom[1821] = 8'hd3 ;
            rom[1822] = 8'h08 ;
            rom[1823] = 8'he9 ;
            rom[1824] = 8'hbd ;
            rom[1825] = 8'h1b ;
            rom[1826] = 8'hd7 ;
            rom[1827] = 8'he0 ;
            rom[1828] = 8'hdd ;
            rom[1829] = 8'hf7 ;
            rom[1830] = 8'h03 ;
            rom[1831] = 8'h15 ;
            rom[1832] = 8'he9 ;
            rom[1833] = 8'hf6 ;
            rom[1834] = 8'hd6 ;
            rom[1835] = 8'hf2 ;
            rom[1836] = 8'hf9 ;
            rom[1837] = 8'he2 ;
            rom[1838] = 8'hfa ;
            rom[1839] = 8'hc0 ;
            rom[1840] = 8'hec ;
            rom[1841] = 8'h08 ;
            rom[1842] = 8'hdf ;
            rom[1843] = 8'h03 ;
            rom[1844] = 8'h0e ;
            rom[1845] = 8'h03 ;
            rom[1846] = 8'hd5 ;
            rom[1847] = 8'hce ;
            rom[1848] = 8'h27 ;
            rom[1849] = 8'hf4 ;
            rom[1850] = 8'h07 ;
            rom[1851] = 8'hd4 ;
            rom[1852] = 8'h01 ;
            rom[1853] = 8'hd5 ;
            rom[1854] = 8'h03 ;
            rom[1855] = 8'h10 ;
            rom[1856] = 8'hde ;
            rom[1857] = 8'hfa ;
            rom[1858] = 8'hf7 ;
            rom[1859] = 8'heb ;
            rom[1860] = 8'hfe ;
            rom[1861] = 8'hbb ;
            rom[1862] = 8'he3 ;
            rom[1863] = 8'hf6 ;
            rom[1864] = 8'h06 ;
            rom[1865] = 8'hf1 ;
            rom[1866] = 8'h1c ;
            rom[1867] = 8'hec ;
            rom[1868] = 8'hf8 ;
            rom[1869] = 8'h0d ;
            rom[1870] = 8'he4 ;
            rom[1871] = 8'h26 ;
            rom[1872] = 8'he8 ;
            rom[1873] = 8'h03 ;
            rom[1874] = 8'hf0 ;
            rom[1875] = 8'h0c ;
            rom[1876] = 8'h04 ;
            rom[1877] = 8'hf5 ;
            rom[1878] = 8'hf2 ;
            rom[1879] = 8'he9 ;
            rom[1880] = 8'h2a ;
            rom[1881] = 8'h02 ;
            rom[1882] = 8'h11 ;
            rom[1883] = 8'h1c ;
            rom[1884] = 8'h1d ;
            rom[1885] = 8'h01 ;
            rom[1886] = 8'hf0 ;
            rom[1887] = 8'hec ;
            rom[1888] = 8'h0b ;
            rom[1889] = 8'hde ;
            rom[1890] = 8'h25 ;
            rom[1891] = 8'he9 ;
            rom[1892] = 8'h23 ;
            rom[1893] = 8'hde ;
            rom[1894] = 8'h19 ;
            rom[1895] = 8'h08 ;
            rom[1896] = 8'hda ;
            rom[1897] = 8'h0d ;
            rom[1898] = 8'hfc ;
            rom[1899] = 8'hd8 ;
            rom[1900] = 8'he6 ;
            rom[1901] = 8'h08 ;
            rom[1902] = 8'h02 ;
            rom[1903] = 8'h0d ;
            rom[1904] = 8'h26 ;
            rom[1905] = 8'hf0 ;
            rom[1906] = 8'h09 ;
            rom[1907] = 8'hfc ;
            rom[1908] = 8'hf0 ;
            rom[1909] = 8'hd8 ;
            rom[1910] = 8'hef ;
            rom[1911] = 8'h20 ;
            rom[1912] = 8'h11 ;
            rom[1913] = 8'h19 ;
            rom[1914] = 8'h1d ;
            rom[1915] = 8'hd8 ;
            rom[1916] = 8'hf5 ;
            rom[1917] = 8'hf1 ;
            rom[1918] = 8'hc7 ;
            rom[1919] = 8'hcd ;
            rom[1920] = 8'he9 ;
            rom[1921] = 8'hd9 ;
            rom[1922] = 8'h03 ;
            rom[1923] = 8'h3a ;
            rom[1924] = 8'hfc ;
            rom[1925] = 8'hff ;
            rom[1926] = 8'h00 ;
            rom[1927] = 8'hfa ;
            rom[1928] = 8'he4 ;
            rom[1929] = 8'h0f ;
            rom[1930] = 8'hc9 ;
            rom[1931] = 8'hd6 ;
            rom[1932] = 8'hd7 ;
            rom[1933] = 8'h0d ;
            rom[1934] = 8'h10 ;
            rom[1935] = 8'h11 ;
            rom[1936] = 8'hf0 ;
            rom[1937] = 8'h29 ;
            rom[1938] = 8'he3 ;
            rom[1939] = 8'h00 ;
            rom[1940] = 8'h14 ;
            rom[1941] = 8'h07 ;
            rom[1942] = 8'hfc ;
            rom[1943] = 8'h16 ;
            rom[1944] = 8'h14 ;
            rom[1945] = 8'h11 ;
            rom[1946] = 8'h0d ;
            rom[1947] = 8'h16 ;
            rom[1948] = 8'h08 ;
            rom[1949] = 8'hfa ;
            rom[1950] = 8'hec ;
            rom[1951] = 8'hfb ;
            rom[1952] = 8'h26 ;
            rom[1953] = 8'hf8 ;
            rom[1954] = 8'hdb ;
            rom[1955] = 8'hf7 ;
            rom[1956] = 8'heb ;
            rom[1957] = 8'hef ;
            rom[1958] = 8'h0f ;
            rom[1959] = 8'he7 ;
            rom[1960] = 8'h14 ;
            rom[1961] = 8'h00 ;
            rom[1962] = 8'hf6 ;
            rom[1963] = 8'h0d ;
            rom[1964] = 8'h0d ;
            rom[1965] = 8'h02 ;
            rom[1966] = 8'hf6 ;
            rom[1967] = 8'h0e ;
            rom[1968] = 8'hf6 ;
            rom[1969] = 8'h14 ;
            rom[1970] = 8'hf2 ;
            rom[1971] = 8'h18 ;
            rom[1972] = 8'hff ;
            rom[1973] = 8'h0b ;
            rom[1974] = 8'hc5 ;
            rom[1975] = 8'heb ;
            rom[1976] = 8'hea ;
            rom[1977] = 8'h04 ;
            rom[1978] = 8'h23 ;
            rom[1979] = 8'h19 ;
            rom[1980] = 8'hf2 ;
            rom[1981] = 8'h0d ;
            rom[1982] = 8'hea ;
            rom[1983] = 8'h03 ;
            rom[1984] = 8'hfb ;
            rom[1985] = 8'h0a ;
            rom[1986] = 8'h0f ;
            rom[1987] = 8'heb ;
            rom[1988] = 8'hfc ;
            rom[1989] = 8'hd2 ;
            rom[1990] = 8'hf0 ;
            rom[1991] = 8'hff ;
            rom[1992] = 8'h0c ;
            rom[1993] = 8'hed ;
            rom[1994] = 8'h13 ;
            rom[1995] = 8'h17 ;
            rom[1996] = 8'h0c ;
            rom[1997] = 8'h0b ;
            rom[1998] = 8'hdf ;
            rom[1999] = 8'hdf ;
            rom[2000] = 8'h08 ;
            rom[2001] = 8'h23 ;
            rom[2002] = 8'hdc ;
            rom[2003] = 8'hfa ;
            rom[2004] = 8'he6 ;
            rom[2005] = 8'h02 ;
            rom[2006] = 8'h03 ;
            rom[2007] = 8'he0 ;
            rom[2008] = 8'h36 ;
            rom[2009] = 8'hda ;
            rom[2010] = 8'h1a ;
            rom[2011] = 8'h0c ;
            rom[2012] = 8'h08 ;
            rom[2013] = 8'h06 ;
            rom[2014] = 8'h01 ;
            rom[2015] = 8'he7 ;
            rom[2016] = 8'heb ;
            rom[2017] = 8'h27 ;
            rom[2018] = 8'he9 ;
            rom[2019] = 8'he7 ;
            rom[2020] = 8'h12 ;
            rom[2021] = 8'hdb ;
            rom[2022] = 8'hfe ;
            rom[2023] = 8'he3 ;
            rom[2024] = 8'hf3 ;
            rom[2025] = 8'h11 ;
            rom[2026] = 8'hf7 ;
            rom[2027] = 8'hf8 ;
            rom[2028] = 8'he5 ;
            rom[2029] = 8'hf0 ;
            rom[2030] = 8'hf7 ;
            rom[2031] = 8'hf1 ;
            rom[2032] = 8'h17 ;
            rom[2033] = 8'h19 ;
            rom[2034] = 8'hf3 ;
            rom[2035] = 8'hf4 ;
            rom[2036] = 8'h0e ;
            rom[2037] = 8'he3 ;
            rom[2038] = 8'hfc ;
            rom[2039] = 8'hf8 ;
            rom[2040] = 8'hfb ;
            rom[2041] = 8'he8 ;
            rom[2042] = 8'h08 ;
            rom[2043] = 8'h03 ;
            rom[2044] = 8'hf7 ;
            rom[2045] = 8'hdd ;
            rom[2046] = 8'hfd ;
            rom[2047] = 8'he8 ;
            rom[2048] = 8'hf5 ;
            rom[2049] = 8'he5 ;
            rom[2050] = 8'hfc ;
            rom[2051] = 8'h1d ;
            rom[2052] = 8'h10 ;
            rom[2053] = 8'h02 ;
            rom[2054] = 8'h0c ;
            rom[2055] = 8'h2e ;
            rom[2056] = 8'heb ;
            rom[2057] = 8'hfe ;
            rom[2058] = 8'he5 ;
            rom[2059] = 8'hcb ;
            rom[2060] = 8'hf1 ;
            rom[2061] = 8'h0a ;
            rom[2062] = 8'h16 ;
            rom[2063] = 8'hf9 ;
            rom[2064] = 8'hfc ;
            rom[2065] = 8'hfa ;
            rom[2066] = 8'he8 ;
            rom[2067] = 8'h02 ;
            rom[2068] = 8'he0 ;
            rom[2069] = 8'hef ;
            rom[2070] = 8'hfd ;
            rom[2071] = 8'he3 ;
            rom[2072] = 8'hf1 ;
            rom[2073] = 8'h04 ;
            rom[2074] = 8'h1b ;
            rom[2075] = 8'hf5 ;
            rom[2076] = 8'h18 ;
            rom[2077] = 8'he9 ;
            rom[2078] = 8'hd8 ;
            rom[2079] = 8'hfc ;
            rom[2080] = 8'h1b ;
            rom[2081] = 8'h1a ;
            rom[2082] = 8'hcd ;
            rom[2083] = 8'h13 ;
            rom[2084] = 8'he8 ;
            rom[2085] = 8'h01 ;
            rom[2086] = 8'h37 ;
            rom[2087] = 8'hf9 ;
            rom[2088] = 8'h04 ;
            rom[2089] = 8'h0d ;
            rom[2090] = 8'h0a ;
            rom[2091] = 8'h08 ;
            rom[2092] = 8'h11 ;
            rom[2093] = 8'hee ;
            rom[2094] = 8'h12 ;
            rom[2095] = 8'h19 ;
            rom[2096] = 8'h02 ;
            rom[2097] = 8'h1a ;
            rom[2098] = 8'h12 ;
            rom[2099] = 8'h00 ;
            rom[2100] = 8'hf4 ;
            rom[2101] = 8'h0e ;
            rom[2102] = 8'h15 ;
            rom[2103] = 8'hc5 ;
            rom[2104] = 8'hed ;
            rom[2105] = 8'hf4 ;
            rom[2106] = 8'h16 ;
            rom[2107] = 8'hfe ;
            rom[2108] = 8'hf8 ;
            rom[2109] = 8'h04 ;
            rom[2110] = 8'hea ;
            rom[2111] = 8'h09 ;
            rom[2112] = 8'h25 ;
            rom[2113] = 8'h0a ;
            rom[2114] = 8'h01 ;
            rom[2115] = 8'hde ;
            rom[2116] = 8'hdf ;
            rom[2117] = 8'he6 ;
            rom[2118] = 8'heb ;
            rom[2119] = 8'h15 ;
            rom[2120] = 8'h24 ;
            rom[2121] = 8'hf8 ;
            rom[2122] = 8'hde ;
            rom[2123] = 8'h1c ;
            rom[2124] = 8'hf9 ;
            rom[2125] = 8'h0b ;
            rom[2126] = 8'h21 ;
            rom[2127] = 8'h21 ;
            rom[2128] = 8'h18 ;
            rom[2129] = 8'hec ;
            rom[2130] = 8'hdd ;
            rom[2131] = 8'he3 ;
            rom[2132] = 8'h00 ;
            rom[2133] = 8'he0 ;
            rom[2134] = 8'hfe ;
            rom[2135] = 8'h10 ;
            rom[2136] = 8'h0c ;
            rom[2137] = 8'hfd ;
            rom[2138] = 8'h06 ;
            rom[2139] = 8'hce ;
            rom[2140] = 8'heb ;
            rom[2141] = 8'hee ;
            rom[2142] = 8'h06 ;
            rom[2143] = 8'h1b ;
            rom[2144] = 8'he2 ;
            rom[2145] = 8'h1c ;
            rom[2146] = 8'hf2 ;
            rom[2147] = 8'hba ;
            rom[2148] = 8'h16 ;
            rom[2149] = 8'hce ;
            rom[2150] = 8'hff ;
            rom[2151] = 8'h36 ;
            rom[2152] = 8'hfe ;
            rom[2153] = 8'h19 ;
            rom[2154] = 8'h05 ;
            rom[2155] = 8'hee ;
            rom[2156] = 8'hea ;
            rom[2157] = 8'h0e ;
            rom[2158] = 8'hf4 ;
            rom[2159] = 8'h18 ;
            rom[2160] = 8'h0c ;
            rom[2161] = 8'h19 ;
            rom[2162] = 8'h37 ;
            rom[2163] = 8'h0d ;
            rom[2164] = 8'heb ;
            rom[2165] = 8'hea ;
            rom[2166] = 8'h08 ;
            rom[2167] = 8'h1f ;
            rom[2168] = 8'h01 ;
            rom[2169] = 8'h1b ;
            rom[2170] = 8'h13 ;
            rom[2171] = 8'hf5 ;
            rom[2172] = 8'hfe ;
            rom[2173] = 8'hfb ;
            rom[2174] = 8'he6 ;
            rom[2175] = 8'h11 ;
            rom[2176] = 8'h00 ;
            rom[2177] = 8'he4 ;
            rom[2178] = 8'h08 ;
            rom[2179] = 8'h03 ;
            rom[2180] = 8'hfe ;
            rom[2181] = 8'hdf ;
            rom[2182] = 8'h10 ;
            rom[2183] = 8'h28 ;
            rom[2184] = 8'hda ;
            rom[2185] = 8'heb ;
            rom[2186] = 8'hf1 ;
            rom[2187] = 8'hdd ;
            rom[2188] = 8'hfe ;
            rom[2189] = 8'hd6 ;
            rom[2190] = 8'hf8 ;
            rom[2191] = 8'hd9 ;
            rom[2192] = 8'he9 ;
            rom[2193] = 8'he0 ;
            rom[2194] = 8'h0c ;
            rom[2195] = 8'h00 ;
            rom[2196] = 8'h05 ;
            rom[2197] = 8'hfc ;
            rom[2198] = 8'h09 ;
            rom[2199] = 8'hf4 ;
            rom[2200] = 8'hd0 ;
            rom[2201] = 8'h0b ;
            rom[2202] = 8'h11 ;
            rom[2203] = 8'he2 ;
            rom[2204] = 8'h0a ;
            rom[2205] = 8'he4 ;
            rom[2206] = 8'h15 ;
            rom[2207] = 8'h17 ;
            rom[2208] = 8'h21 ;
            rom[2209] = 8'hff ;
            rom[2210] = 8'hfb ;
            rom[2211] = 8'hda ;
            rom[2212] = 8'he5 ;
            rom[2213] = 8'h15 ;
            rom[2214] = 8'hfb ;
            rom[2215] = 8'hf0 ;
            rom[2216] = 8'hf8 ;
            rom[2217] = 8'he6 ;
            rom[2218] = 8'hf6 ;
            rom[2219] = 8'hd7 ;
            rom[2220] = 8'h01 ;
            rom[2221] = 8'h1f ;
            rom[2222] = 8'he1 ;
            rom[2223] = 8'h0a ;
            rom[2224] = 8'h03 ;
            rom[2225] = 8'heb ;
            rom[2226] = 8'hea ;
            rom[2227] = 8'h11 ;
            rom[2228] = 8'hf1 ;
            rom[2229] = 8'hfd ;
            rom[2230] = 8'h19 ;
            rom[2231] = 8'hfd ;
            rom[2232] = 8'hdd ;
            rom[2233] = 8'hfd ;
            rom[2234] = 8'h22 ;
            rom[2235] = 8'h0b ;
            rom[2236] = 8'h12 ;
            rom[2237] = 8'h28 ;
            rom[2238] = 8'hd7 ;
            rom[2239] = 8'h03 ;
            rom[2240] = 8'hf4 ;
            rom[2241] = 8'h12 ;
            rom[2242] = 8'he6 ;
            rom[2243] = 8'hfc ;
            rom[2244] = 8'hee ;
            rom[2245] = 8'hf1 ;
            rom[2246] = 8'h16 ;
            rom[2247] = 8'h0d ;
            rom[2248] = 8'hf7 ;
            rom[2249] = 8'hea ;
            rom[2250] = 8'hd6 ;
            rom[2251] = 8'h08 ;
            rom[2252] = 8'h15 ;
            rom[2253] = 8'he6 ;
            rom[2254] = 8'h02 ;
            rom[2255] = 8'h02 ;
            rom[2256] = 8'h13 ;
            rom[2257] = 8'hfc ;
            rom[2258] = 8'h13 ;
            rom[2259] = 8'hde ;
            rom[2260] = 8'he8 ;
            rom[2261] = 8'he8 ;
            rom[2262] = 8'h1d ;
            rom[2263] = 8'hff ;
            rom[2264] = 8'h02 ;
            rom[2265] = 8'h05 ;
            rom[2266] = 8'h34 ;
            rom[2267] = 8'h0f ;
            rom[2268] = 8'hf3 ;
            rom[2269] = 8'hdc ;
            rom[2270] = 8'hfe ;
            rom[2271] = 8'he5 ;
            rom[2272] = 8'hf3 ;
            rom[2273] = 8'h00 ;
            rom[2274] = 8'hec ;
            rom[2275] = 8'hff ;
            rom[2276] = 8'h08 ;
            rom[2277] = 8'h18 ;
            rom[2278] = 8'h00 ;
            rom[2279] = 8'hfe ;
            rom[2280] = 8'h02 ;
            rom[2281] = 8'h00 ;
            rom[2282] = 8'h39 ;
            rom[2283] = 8'h16 ;
            rom[2284] = 8'hfd ;
            rom[2285] = 8'h14 ;
            rom[2286] = 8'he3 ;
            rom[2287] = 8'hf0 ;
            rom[2288] = 8'h08 ;
            rom[2289] = 8'heb ;
            rom[2290] = 8'h1a ;
            rom[2291] = 8'he4 ;
            rom[2292] = 8'he4 ;
            rom[2293] = 8'h13 ;
            rom[2294] = 8'he5 ;
            rom[2295] = 8'h04 ;
            rom[2296] = 8'h0f ;
            rom[2297] = 8'h26 ;
            rom[2298] = 8'hf3 ;
            rom[2299] = 8'h02 ;
            rom[2300] = 8'hf0 ;
            rom[2301] = 8'hf3 ;
            rom[2302] = 8'heb ;
            rom[2303] = 8'hc1 ;
            rom[2304] = 8'h16 ;
            rom[2305] = 8'hd7 ;
            rom[2306] = 8'h0e ;
            rom[2307] = 8'h00 ;
            rom[2308] = 8'hf6 ;
            rom[2309] = 8'h17 ;
            rom[2310] = 8'h01 ;
            rom[2311] = 8'hfc ;
            rom[2312] = 8'h14 ;
            rom[2313] = 8'h17 ;
            rom[2314] = 8'h01 ;
            rom[2315] = 8'h11 ;
            rom[2316] = 8'h07 ;
            rom[2317] = 8'hd2 ;
            rom[2318] = 8'h29 ;
            rom[2319] = 8'hfe ;
            rom[2320] = 8'hf3 ;
            rom[2321] = 8'h04 ;
            rom[2322] = 8'hdb ;
            rom[2323] = 8'h04 ;
            rom[2324] = 8'h0d ;
            rom[2325] = 8'hf2 ;
            rom[2326] = 8'h09 ;
            rom[2327] = 8'h01 ;
            rom[2328] = 8'hfc ;
            rom[2329] = 8'hf8 ;
            rom[2330] = 8'h09 ;
            rom[2331] = 8'hf2 ;
            rom[2332] = 8'h05 ;
            rom[2333] = 8'hfa ;
            rom[2334] = 8'h08 ;
            rom[2335] = 8'he0 ;
            rom[2336] = 8'hf0 ;
            rom[2337] = 8'h0a ;
            rom[2338] = 8'hdc ;
            rom[2339] = 8'h06 ;
            rom[2340] = 8'hf8 ;
            rom[2341] = 8'h27 ;
            rom[2342] = 8'hde ;
            rom[2343] = 8'hcb ;
            rom[2344] = 8'h02 ;
            rom[2345] = 8'hf9 ;
            rom[2346] = 8'h17 ;
            rom[2347] = 8'hff ;
            rom[2348] = 8'h31 ;
            rom[2349] = 8'he7 ;
            rom[2350] = 8'h00 ;
            rom[2351] = 8'hea ;
            rom[2352] = 8'he9 ;
            rom[2353] = 8'h11 ;
            rom[2354] = 8'hee ;
            rom[2355] = 8'hf0 ;
            rom[2356] = 8'h24 ;
            rom[2357] = 8'h10 ;
            rom[2358] = 8'hc5 ;
            rom[2359] = 8'heb ;
            rom[2360] = 8'h00 ;
            rom[2361] = 8'h22 ;
            rom[2362] = 8'h02 ;
            rom[2363] = 8'hf4 ;
            rom[2364] = 8'hfa ;
            rom[2365] = 8'hfc ;
            rom[2366] = 8'h02 ;
            rom[2367] = 8'he1 ;
            rom[2368] = 8'he1 ;
            rom[2369] = 8'h03 ;
            rom[2370] = 8'hf8 ;
            rom[2371] = 8'h11 ;
            rom[2372] = 8'hf0 ;
            rom[2373] = 8'h0d ;
            rom[2374] = 8'h02 ;
            rom[2375] = 8'hf5 ;
            rom[2376] = 8'h08 ;
            rom[2377] = 8'h03 ;
            rom[2378] = 8'he5 ;
            rom[2379] = 8'hfa ;
            rom[2380] = 8'heb ;
            rom[2381] = 8'h26 ;
            rom[2382] = 8'hf5 ;
            rom[2383] = 8'h15 ;
            rom[2384] = 8'h2a ;
            rom[2385] = 8'h0c ;
            rom[2386] = 8'h16 ;
            rom[2387] = 8'h02 ;
            rom[2388] = 8'hee ;
            rom[2389] = 8'hdc ;
            rom[2390] = 8'h01 ;
            rom[2391] = 8'hfa ;
            rom[2392] = 8'h04 ;
            rom[2393] = 8'hff ;
            rom[2394] = 8'hdd ;
            rom[2395] = 8'h0e ;
            rom[2396] = 8'h02 ;
            rom[2397] = 8'hcf ;
            rom[2398] = 8'h24 ;
            rom[2399] = 8'h15 ;
            rom[2400] = 8'hf7 ;
            rom[2401] = 8'h37 ;
            rom[2402] = 8'hf9 ;
            rom[2403] = 8'hdc ;
            rom[2404] = 8'hdd ;
            rom[2405] = 8'he8 ;
            rom[2406] = 8'hf1 ;
            rom[2407] = 8'he6 ;
            rom[2408] = 8'h06 ;
            rom[2409] = 8'h04 ;
            rom[2410] = 8'he4 ;
            rom[2411] = 8'hf5 ;
            rom[2412] = 8'h02 ;
            rom[2413] = 8'hda ;
            rom[2414] = 8'h11 ;
            rom[2415] = 8'hda ;
            rom[2416] = 8'h00 ;
            rom[2417] = 8'hdf ;
            rom[2418] = 8'h07 ;
            rom[2419] = 8'hf5 ;
            rom[2420] = 8'hf2 ;
            rom[2421] = 8'h08 ;
            rom[2422] = 8'h26 ;
            rom[2423] = 8'hf4 ;
            rom[2424] = 8'hff ;
            rom[2425] = 8'he8 ;
            rom[2426] = 8'h23 ;
            rom[2427] = 8'hd1 ;
            rom[2428] = 8'h02 ;
            rom[2429] = 8'hcc ;
            rom[2430] = 8'he8 ;
            rom[2431] = 8'he4 ;
            rom[2432] = 8'hee ;
            rom[2433] = 8'hcb ;
            rom[2434] = 8'hd9 ;
            rom[2435] = 8'h0f ;
            rom[2436] = 8'h03 ;
            rom[2437] = 8'h06 ;
            rom[2438] = 8'he8 ;
            rom[2439] = 8'h21 ;
            rom[2440] = 8'h0f ;
            rom[2441] = 8'h05 ;
            rom[2442] = 8'h1f ;
            rom[2443] = 8'hec ;
            rom[2444] = 8'h06 ;
            rom[2445] = 8'h03 ;
            rom[2446] = 8'h0a ;
            rom[2447] = 8'hd5 ;
            rom[2448] = 8'hfa ;
            rom[2449] = 8'h0a ;
            rom[2450] = 8'h01 ;
            rom[2451] = 8'he7 ;
            rom[2452] = 8'h0a ;
            rom[2453] = 8'h06 ;
            rom[2454] = 8'h04 ;
            rom[2455] = 8'hdd ;
            rom[2456] = 8'hf4 ;
            rom[2457] = 8'h19 ;
            rom[2458] = 8'hf5 ;
            rom[2459] = 8'hf7 ;
            rom[2460] = 8'h0b ;
            rom[2461] = 8'h11 ;
            rom[2462] = 8'h03 ;
            rom[2463] = 8'h1c ;
            rom[2464] = 8'h0a ;
            rom[2465] = 8'hdc ;
            rom[2466] = 8'hdb ;
            rom[2467] = 8'h14 ;
            rom[2468] = 8'he0 ;
            rom[2469] = 8'h0e ;
            rom[2470] = 8'h1c ;
            rom[2471] = 8'h15 ;
            rom[2472] = 8'h10 ;
            rom[2473] = 8'h02 ;
            rom[2474] = 8'h0d ;
            rom[2475] = 8'h01 ;
            rom[2476] = 8'h22 ;
            rom[2477] = 8'h09 ;
            rom[2478] = 8'hf5 ;
            rom[2479] = 8'h0d ;
            rom[2480] = 8'he6 ;
            rom[2481] = 8'h01 ;
            rom[2482] = 8'h38 ;
            rom[2483] = 8'h0b ;
            rom[2484] = 8'h09 ;
            rom[2485] = 8'hff ;
            rom[2486] = 8'h21 ;
            rom[2487] = 8'h12 ;
            rom[2488] = 8'hef ;
            rom[2489] = 8'hf4 ;
            rom[2490] = 8'hfd ;
            rom[2491] = 8'hfe ;
            rom[2492] = 8'he5 ;
            rom[2493] = 8'h0b ;
            rom[2494] = 8'he3 ;
            rom[2495] = 8'h1c ;
            rom[2496] = 8'h27 ;
            rom[2497] = 8'h11 ;
            rom[2498] = 8'hf3 ;
            rom[2499] = 8'hfa ;
            rom[2500] = 8'h08 ;
            rom[2501] = 8'h05 ;
            rom[2502] = 8'h14 ;
            rom[2503] = 8'h0f ;
            rom[2504] = 8'h38 ;
            rom[2505] = 8'hd5 ;
            rom[2506] = 8'hc5 ;
            rom[2507] = 8'h0b ;
            rom[2508] = 8'hff ;
            rom[2509] = 8'hee ;
            rom[2510] = 8'h16 ;
            rom[2511] = 8'h05 ;
            rom[2512] = 8'h00 ;
            rom[2513] = 8'h0e ;
            rom[2514] = 8'hfb ;
            rom[2515] = 8'he6 ;
            rom[2516] = 8'he2 ;
            rom[2517] = 8'h1a ;
            rom[2518] = 8'h0c ;
            rom[2519] = 8'hfc ;
            rom[2520] = 8'h05 ;
            rom[2521] = 8'h10 ;
            rom[2522] = 8'h15 ;
            rom[2523] = 8'hf5 ;
            rom[2524] = 8'h17 ;
            rom[2525] = 8'hed ;
            rom[2526] = 8'h19 ;
            rom[2527] = 8'h09 ;
            rom[2528] = 8'hf4 ;
            rom[2529] = 8'h4a ;
            rom[2530] = 8'h09 ;
            rom[2531] = 8'hd4 ;
            rom[2532] = 8'h08 ;
            rom[2533] = 8'hf7 ;
            rom[2534] = 8'h09 ;
            rom[2535] = 8'h1f ;
            rom[2536] = 8'h20 ;
            rom[2537] = 8'h03 ;
            rom[2538] = 8'hfb ;
            rom[2539] = 8'he3 ;
            rom[2540] = 8'h09 ;
            rom[2541] = 8'hfb ;
            rom[2542] = 8'he0 ;
            rom[2543] = 8'h11 ;
            rom[2544] = 8'h05 ;
            rom[2545] = 8'h20 ;
            rom[2546] = 8'h2e ;
            rom[2547] = 8'hf7 ;
            rom[2548] = 8'hea ;
            rom[2549] = 8'hd2 ;
            rom[2550] = 8'h24 ;
            rom[2551] = 8'hfa ;
            rom[2552] = 8'hed ;
            rom[2553] = 8'h0b ;
            rom[2554] = 8'h2b ;
            rom[2555] = 8'he9 ;
            rom[2556] = 8'hec ;
            rom[2557] = 8'h15 ;
            rom[2558] = 8'h04 ;
            rom[2559] = 8'hfa ;
            rom[2560] = 8'h0d ;
            rom[2561] = 8'h12 ;
            rom[2562] = 8'he9 ;
            rom[2563] = 8'h29 ;
            rom[2564] = 8'h21 ;
            rom[2565] = 8'he1 ;
            rom[2566] = 8'he8 ;
            rom[2567] = 8'hf7 ;
            rom[2568] = 8'he6 ;
            rom[2569] = 8'h04 ;
            rom[2570] = 8'he0 ;
            rom[2571] = 8'he8 ;
            rom[2572] = 8'hf4 ;
            rom[2573] = 8'hfb ;
            rom[2574] = 8'hd5 ;
            rom[2575] = 8'h01 ;
            rom[2576] = 8'hf8 ;
            rom[2577] = 8'h2a ;
            rom[2578] = 8'hf2 ;
            rom[2579] = 8'hdc ;
            rom[2580] = 8'h19 ;
            rom[2581] = 8'h0a ;
            rom[2582] = 8'hd6 ;
            rom[2583] = 8'hff ;
            rom[2584] = 8'hf9 ;
            rom[2585] = 8'h0d ;
            rom[2586] = 8'hf8 ;
            rom[2587] = 8'h09 ;
            rom[2588] = 8'h18 ;
            rom[2589] = 8'hfd ;
            rom[2590] = 8'h09 ;
            rom[2591] = 8'h06 ;
            rom[2592] = 8'hd7 ;
            rom[2593] = 8'hf0 ;
            rom[2594] = 8'hf8 ;
            rom[2595] = 8'h23 ;
            rom[2596] = 8'hcc ;
            rom[2597] = 8'h01 ;
            rom[2598] = 8'hf2 ;
            rom[2599] = 8'h17 ;
            rom[2600] = 8'hf3 ;
            rom[2601] = 8'hf0 ;
            rom[2602] = 8'he5 ;
            rom[2603] = 8'hf6 ;
            rom[2604] = 8'h0f ;
            rom[2605] = 8'hf2 ;
            rom[2606] = 8'h09 ;
            rom[2607] = 8'hfb ;
            rom[2608] = 8'hed ;
            rom[2609] = 8'he3 ;
            rom[2610] = 8'he6 ;
            rom[2611] = 8'h04 ;
            rom[2612] = 8'h0a ;
            rom[2613] = 8'hf2 ;
            rom[2614] = 8'he3 ;
            rom[2615] = 8'hf6 ;
            rom[2616] = 8'h25 ;
            rom[2617] = 8'hda ;
            rom[2618] = 8'h03 ;
            rom[2619] = 8'h01 ;
            rom[2620] = 8'hf0 ;
            rom[2621] = 8'he7 ;
            rom[2622] = 8'h1a ;
            rom[2623] = 8'h0e ;
            rom[2624] = 8'h01 ;
            rom[2625] = 8'hec ;
            rom[2626] = 8'hc0 ;
            rom[2627] = 8'hef ;
            rom[2628] = 8'hff ;
            rom[2629] = 8'hc9 ;
            rom[2630] = 8'hf5 ;
            rom[2631] = 8'hf2 ;
            rom[2632] = 8'h05 ;
            rom[2633] = 8'h17 ;
            rom[2634] = 8'h3c ;
            rom[2635] = 8'h2a ;
            rom[2636] = 8'h03 ;
            rom[2637] = 8'h0d ;
            rom[2638] = 8'hfb ;
            rom[2639] = 8'h26 ;
            rom[2640] = 8'hdc ;
            rom[2641] = 8'h1e ;
            rom[2642] = 8'hd8 ;
            rom[2643] = 8'h18 ;
            rom[2644] = 8'h05 ;
            rom[2645] = 8'h02 ;
            rom[2646] = 8'h02 ;
            rom[2647] = 8'hf3 ;
            rom[2648] = 8'hf5 ;
            rom[2649] = 8'h0d ;
            rom[2650] = 8'he3 ;
            rom[2651] = 8'h0d ;
            rom[2652] = 8'h10 ;
            rom[2653] = 8'h0e ;
            rom[2654] = 8'h0a ;
            rom[2655] = 8'h04 ;
            rom[2656] = 8'he7 ;
            rom[2657] = 8'ha8 ;
            rom[2658] = 8'hf5 ;
            rom[2659] = 8'he8 ;
            rom[2660] = 8'hfd ;
            rom[2661] = 8'hce ;
            rom[2662] = 8'hfd ;
            rom[2663] = 8'h06 ;
            rom[2664] = 8'hc9 ;
            rom[2665] = 8'hf8 ;
            rom[2666] = 8'hbc ;
            rom[2667] = 8'he0 ;
            rom[2668] = 8'hf3 ;
            rom[2669] = 8'hd6 ;
            rom[2670] = 8'hf4 ;
            rom[2671] = 8'h01 ;
            rom[2672] = 8'hf2 ;
            rom[2673] = 8'hef ;
            rom[2674] = 8'hfd ;
            rom[2675] = 8'h06 ;
            rom[2676] = 8'h1c ;
            rom[2677] = 8'h10 ;
            rom[2678] = 8'hf9 ;
            rom[2679] = 8'h01 ;
            rom[2680] = 8'hf6 ;
            rom[2681] = 8'h1b ;
            rom[2682] = 8'hde ;
            rom[2683] = 8'h2d ;
            rom[2684] = 8'hfc ;
            rom[2685] = 8'h02 ;
            rom[2686] = 8'hee ;
            rom[2687] = 8'h00 ;
            rom[2688] = 8'hd6 ;
            rom[2689] = 8'hf5 ;
            rom[2690] = 8'hf4 ;
            rom[2691] = 8'hfb ;
            rom[2692] = 8'hfb ;
            rom[2693] = 8'hb4 ;
            rom[2694] = 8'hf9 ;
            rom[2695] = 8'hfa ;
            rom[2696] = 8'he8 ;
            rom[2697] = 8'hfa ;
            rom[2698] = 8'he1 ;
            rom[2699] = 8'hf2 ;
            rom[2700] = 8'hc8 ;
            rom[2701] = 8'h27 ;
            rom[2702] = 8'hed ;
            rom[2703] = 8'h1b ;
            rom[2704] = 8'h2e ;
            rom[2705] = 8'hdf ;
            rom[2706] = 8'h08 ;
            rom[2707] = 8'hdb ;
            rom[2708] = 8'hfd ;
            rom[2709] = 8'he7 ;
            rom[2710] = 8'h12 ;
            rom[2711] = 8'h0e ;
            rom[2712] = 8'he3 ;
            rom[2713] = 8'h06 ;
            rom[2714] = 8'h15 ;
            rom[2715] = 8'hfd ;
            rom[2716] = 8'hf3 ;
            rom[2717] = 8'h1a ;
            rom[2718] = 8'hf6 ;
            rom[2719] = 8'h0c ;
            rom[2720] = 8'hfd ;
            rom[2721] = 8'he4 ;
            rom[2722] = 8'h09 ;
            rom[2723] = 8'hdb ;
            rom[2724] = 8'h12 ;
            rom[2725] = 8'hef ;
            rom[2726] = 8'hfb ;
            rom[2727] = 8'h14 ;
            rom[2728] = 8'h13 ;
            rom[2729] = 8'h16 ;
            rom[2730] = 8'h03 ;
            rom[2731] = 8'hee ;
            rom[2732] = 8'h00 ;
            rom[2733] = 8'h2b ;
            rom[2734] = 8'hdd ;
            rom[2735] = 8'h06 ;
            rom[2736] = 8'h0d ;
            rom[2737] = 8'h38 ;
            rom[2738] = 8'h13 ;
            rom[2739] = 8'h10 ;
            rom[2740] = 8'h21 ;
            rom[2741] = 8'he4 ;
            rom[2742] = 8'hca ;
            rom[2743] = 8'hf7 ;
            rom[2744] = 8'h06 ;
            rom[2745] = 8'h05 ;
            rom[2746] = 8'h22 ;
            rom[2747] = 8'h09 ;
            rom[2748] = 8'he6 ;
            rom[2749] = 8'heb ;
            rom[2750] = 8'h05 ;
            rom[2751] = 8'h02 ;
            rom[2752] = 8'h18 ;
            rom[2753] = 8'h14 ;
            rom[2754] = 8'h0c ;
            rom[2755] = 8'hc4 ;
            rom[2756] = 8'h07 ;
            rom[2757] = 8'hfd ;
            rom[2758] = 8'hef ;
            rom[2759] = 8'hf6 ;
            rom[2760] = 8'he2 ;
            rom[2761] = 8'hdd ;
            rom[2762] = 8'h05 ;
            rom[2763] = 8'h25 ;
            rom[2764] = 8'hfb ;
            rom[2765] = 8'hed ;
            rom[2766] = 8'hfc ;
            rom[2767] = 8'h07 ;
            rom[2768] = 8'hda ;
            rom[2769] = 8'h04 ;
            rom[2770] = 8'h07 ;
            rom[2771] = 8'h05 ;
            rom[2772] = 8'h12 ;
            rom[2773] = 8'hf0 ;
            rom[2774] = 8'hf9 ;
            rom[2775] = 8'hfe ;
            rom[2776] = 8'h34 ;
            rom[2777] = 8'h04 ;
            rom[2778] = 8'h03 ;
            rom[2779] = 8'h03 ;
            rom[2780] = 8'hdb ;
            rom[2781] = 8'h0c ;
            rom[2782] = 8'hd7 ;
            rom[2783] = 8'hea ;
            rom[2784] = 8'h0d ;
            rom[2785] = 8'h09 ;
            rom[2786] = 8'hf7 ;
            rom[2787] = 8'h00 ;
            rom[2788] = 8'h3b ;
            rom[2789] = 8'hfd ;
            rom[2790] = 8'he3 ;
            rom[2791] = 8'he7 ;
            rom[2792] = 8'hea ;
            rom[2793] = 8'h12 ;
            rom[2794] = 8'hfa ;
            rom[2795] = 8'hf4 ;
            rom[2796] = 8'ha7 ;
            rom[2797] = 8'hed ;
            rom[2798] = 8'h04 ;
            rom[2799] = 8'h11 ;
            rom[2800] = 8'he5 ;
            rom[2801] = 8'h14 ;
            rom[2802] = 8'hf8 ;
            rom[2803] = 8'h32 ;
            rom[2804] = 8'h04 ;
            rom[2805] = 8'hdf ;
            rom[2806] = 8'he9 ;
            rom[2807] = 8'h28 ;
            rom[2808] = 8'h0d ;
            rom[2809] = 8'hde ;
            rom[2810] = 8'h04 ;
            rom[2811] = 8'hee ;
            rom[2812] = 8'hd7 ;
            rom[2813] = 8'hdb ;
            rom[2814] = 8'hca ;
            rom[2815] = 8'h20 ;
            rom[2816] = 8'h20 ;
            rom[2817] = 8'h0f ;
            rom[2818] = 8'he5 ;
            rom[2819] = 8'h0d ;
            rom[2820] = 8'he7 ;
            rom[2821] = 8'hc7 ;
            rom[2822] = 8'hed ;
            rom[2823] = 8'hf5 ;
            rom[2824] = 8'h0f ;
            rom[2825] = 8'h35 ;
            rom[2826] = 8'hf4 ;
            rom[2827] = 8'h15 ;
            rom[2828] = 8'he5 ;
            rom[2829] = 8'hff ;
            rom[2830] = 8'hec ;
            rom[2831] = 8'h05 ;
            rom[2832] = 8'hdf ;
            rom[2833] = 8'heb ;
            rom[2834] = 8'hc6 ;
            rom[2835] = 8'h09 ;
            rom[2836] = 8'h0f ;
            rom[2837] = 8'h01 ;
            rom[2838] = 8'h21 ;
            rom[2839] = 8'h08 ;
            rom[2840] = 8'h05 ;
            rom[2841] = 8'hf7 ;
            rom[2842] = 8'hee ;
            rom[2843] = 8'h0b ;
            rom[2844] = 8'h03 ;
            rom[2845] = 8'hf7 ;
            rom[2846] = 8'h20 ;
            rom[2847] = 8'hcf ;
            rom[2848] = 8'hf0 ;
            rom[2849] = 8'h22 ;
            rom[2850] = 8'hee ;
            rom[2851] = 8'he3 ;
            rom[2852] = 8'h09 ;
            rom[2853] = 8'hed ;
            rom[2854] = 8'hbe ;
            rom[2855] = 8'h03 ;
            rom[2856] = 8'hd4 ;
            rom[2857] = 8'he8 ;
            rom[2858] = 8'h10 ;
            rom[2859] = 8'hec ;
            rom[2860] = 8'hdf ;
            rom[2861] = 8'hbe ;
            rom[2862] = 8'he2 ;
            rom[2863] = 8'h1b ;
            rom[2864] = 8'hfa ;
            rom[2865] = 8'h17 ;
            rom[2866] = 8'hf8 ;
            rom[2867] = 8'hce ;
            rom[2868] = 8'hed ;
            rom[2869] = 8'hfa ;
            rom[2870] = 8'hd0 ;
            rom[2871] = 8'he6 ;
            rom[2872] = 8'h2c ;
            rom[2873] = 8'hf9 ;
            rom[2874] = 8'he5 ;
            rom[2875] = 8'he3 ;
            rom[2876] = 8'h16 ;
            rom[2877] = 8'hfa ;
            rom[2878] = 8'hef ;
            rom[2879] = 8'hcc ;
            rom[2880] = 8'hfe ;
            rom[2881] = 8'he3 ;
            rom[2882] = 8'h1a ;
            rom[2883] = 8'he8 ;
            rom[2884] = 8'h14 ;
            rom[2885] = 8'h19 ;
            rom[2886] = 8'hb9 ;
            rom[2887] = 8'hd0 ;
            rom[2888] = 8'he8 ;
            rom[2889] = 8'h02 ;
            rom[2890] = 8'he7 ;
            rom[2891] = 8'hd9 ;
            rom[2892] = 8'h0e ;
            rom[2893] = 8'h0a ;
            rom[2894] = 8'h08 ;
            rom[2895] = 8'h05 ;
            rom[2896] = 8'h12 ;
            rom[2897] = 8'h07 ;
            rom[2898] = 8'h02 ;
            rom[2899] = 8'hf6 ;
            rom[2900] = 8'hf0 ;
            rom[2901] = 8'hc8 ;
            rom[2902] = 8'heb ;
            rom[2903] = 8'hd7 ;
            rom[2904] = 8'h07 ;
            rom[2905] = 8'hd6 ;
            rom[2906] = 8'hda ;
            rom[2907] = 8'hfa ;
            rom[2908] = 8'hd0 ;
            rom[2909] = 8'h10 ;
            rom[2910] = 8'h1e ;
            rom[2911] = 8'hc7 ;
            rom[2912] = 8'h0a ;
            rom[2913] = 8'hf4 ;
            rom[2914] = 8'he8 ;
            rom[2915] = 8'h0e ;
            rom[2916] = 8'h01 ;
            rom[2917] = 8'h09 ;
            rom[2918] = 8'he0 ;
            rom[2919] = 8'h1a ;
            rom[2920] = 8'hc1 ;
            rom[2921] = 8'h09 ;
            rom[2922] = 8'he6 ;
            rom[2923] = 8'he2 ;
            rom[2924] = 8'h07 ;
            rom[2925] = 8'h0c ;
            rom[2926] = 8'hf4 ;
            rom[2927] = 8'hf3 ;
            rom[2928] = 8'hfe ;
            rom[2929] = 8'h1b ;
            rom[2930] = 8'hec ;
            rom[2931] = 8'hf8 ;
            rom[2932] = 8'hd3 ;
            rom[2933] = 8'h08 ;
            rom[2934] = 8'hfc ;
            rom[2935] = 8'hf5 ;
            rom[2936] = 8'h03 ;
            rom[2937] = 8'hf6 ;
            rom[2938] = 8'hd2 ;
            rom[2939] = 8'h1b ;
            rom[2940] = 8'hf5 ;
            rom[2941] = 8'hfa ;
            rom[2942] = 8'h0d ;
            rom[2943] = 8'hf3 ;
            rom[2944] = 8'hda ;
            rom[2945] = 8'hef ;
            rom[2946] = 8'hfc ;
            rom[2947] = 8'hfd ;
            rom[2948] = 8'hbe ;
            rom[2949] = 8'hde ;
            rom[2950] = 8'h15 ;
            rom[2951] = 8'h0e ;
            rom[2952] = 8'hd3 ;
            rom[2953] = 8'h16 ;
            rom[2954] = 8'hcf ;
            rom[2955] = 8'hda ;
            rom[2956] = 8'h06 ;
            rom[2957] = 8'h06 ;
            rom[2958] = 8'h15 ;
            rom[2959] = 8'he2 ;
            rom[2960] = 8'hf5 ;
            rom[2961] = 8'h00 ;
            rom[2962] = 8'hfb ;
            rom[2963] = 8'h0f ;
            rom[2964] = 8'h0e ;
            rom[2965] = 8'he3 ;
            rom[2966] = 8'h07 ;
            rom[2967] = 8'hf4 ;
            rom[2968] = 8'hf6 ;
            rom[2969] = 8'h0d ;
            rom[2970] = 8'h01 ;
            rom[2971] = 8'hd8 ;
            rom[2972] = 8'h00 ;
            rom[2973] = 8'h16 ;
            rom[2974] = 8'hde ;
            rom[2975] = 8'hfc ;
            rom[2976] = 8'h07 ;
            rom[2977] = 8'hd7 ;
            rom[2978] = 8'hff ;
            rom[2979] = 8'hea ;
            rom[2980] = 8'hf7 ;
            rom[2981] = 8'h14 ;
            rom[2982] = 8'h00 ;
            rom[2983] = 8'hd6 ;
            rom[2984] = 8'hfe ;
            rom[2985] = 8'hd4 ;
            rom[2986] = 8'h06 ;
            rom[2987] = 8'he9 ;
            rom[2988] = 8'h24 ;
            rom[2989] = 8'hf4 ;
            rom[2990] = 8'hd6 ;
            rom[2991] = 8'h0a ;
            rom[2992] = 8'h06 ;
            rom[2993] = 8'he7 ;
            rom[2994] = 8'h06 ;
            rom[2995] = 8'h2b ;
            rom[2996] = 8'hfd ;
            rom[2997] = 8'h0e ;
            rom[2998] = 8'hf7 ;
            rom[2999] = 8'hd3 ;
            rom[3000] = 8'he7 ;
            rom[3001] = 8'h27 ;
            rom[3002] = 8'hfe ;
            rom[3003] = 8'h02 ;
            rom[3004] = 8'hdf ;
            rom[3005] = 8'hf4 ;
            rom[3006] = 8'hfa ;
            rom[3007] = 8'h17 ;
            rom[3008] = 8'hfb ;
            rom[3009] = 8'h0a ;
            rom[3010] = 8'hff ;
            rom[3011] = 8'h00 ;
            rom[3012] = 8'h0d ;
            rom[3013] = 8'hea ;
            rom[3014] = 8'he1 ;
            rom[3015] = 8'hed ;
            rom[3016] = 8'hd4 ;
            rom[3017] = 8'h09 ;
            rom[3018] = 8'h10 ;
            rom[3019] = 8'h27 ;
            rom[3020] = 8'hf0 ;
            rom[3021] = 8'h07 ;
            rom[3022] = 8'hf9 ;
            rom[3023] = 8'h00 ;
            rom[3024] = 8'hfb ;
            rom[3025] = 8'h08 ;
            rom[3026] = 8'h05 ;
            rom[3027] = 8'hd0 ;
            rom[3028] = 8'h09 ;
            rom[3029] = 8'hfe ;
            rom[3030] = 8'hfd ;
            rom[3031] = 8'he0 ;
            rom[3032] = 8'hf0 ;
            rom[3033] = 8'he1 ;
            rom[3034] = 8'h17 ;
            rom[3035] = 8'h02 ;
            rom[3036] = 8'h39 ;
            rom[3037] = 8'hfd ;
            rom[3038] = 8'h08 ;
            rom[3039] = 8'he6 ;
            rom[3040] = 8'hfc ;
            rom[3041] = 8'h1c ;
            rom[3042] = 8'h1a ;
            rom[3043] = 8'hff ;
            rom[3044] = 8'he9 ;
            rom[3045] = 8'h0b ;
            rom[3046] = 8'hfa ;
            rom[3047] = 8'hfb ;
            rom[3048] = 8'h01 ;
            rom[3049] = 8'h28 ;
            rom[3050] = 8'h0c ;
            rom[3051] = 8'h03 ;
            rom[3052] = 8'hf8 ;
            rom[3053] = 8'h3a ;
            rom[3054] = 8'hdf ;
            rom[3055] = 8'hfe ;
            rom[3056] = 8'h15 ;
            rom[3057] = 8'h35 ;
            rom[3058] = 8'h17 ;
            rom[3059] = 8'hd8 ;
            rom[3060] = 8'h17 ;
            rom[3061] = 8'hec ;
            rom[3062] = 8'hfa ;
            rom[3063] = 8'h1a ;
            rom[3064] = 8'hfe ;
            rom[3065] = 8'he0 ;
            rom[3066] = 8'h04 ;
            rom[3067] = 8'hed ;
            rom[3068] = 8'h0e ;
            rom[3069] = 8'h0e ;
            rom[3070] = 8'hf6 ;
            rom[3071] = 8'h1f ;
            rom[3072] = 8'hd4 ;
            rom[3073] = 8'hb9 ;
            rom[3074] = 8'hf2 ;
            rom[3075] = 8'he2 ;
            rom[3076] = 8'heb ;
            rom[3077] = 8'h07 ;
            rom[3078] = 8'hf7 ;
            rom[3079] = 8'hfd ;
            rom[3080] = 8'hf2 ;
            rom[3081] = 8'hfe ;
            rom[3082] = 8'h1b ;
            rom[3083] = 8'hf1 ;
            rom[3084] = 8'hfd ;
            rom[3085] = 8'hcc ;
            rom[3086] = 8'h22 ;
            rom[3087] = 8'hfc ;
            rom[3088] = 8'h0c ;
            rom[3089] = 8'heb ;
            rom[3090] = 8'h0f ;
            rom[3091] = 8'h01 ;
            rom[3092] = 8'he8 ;
            rom[3093] = 8'he3 ;
            rom[3094] = 8'hf3 ;
            rom[3095] = 8'hf3 ;
            rom[3096] = 8'h26 ;
            rom[3097] = 8'hf7 ;
            rom[3098] = 8'hf4 ;
            rom[3099] = 8'h14 ;
            rom[3100] = 8'h0c ;
            rom[3101] = 8'h29 ;
            rom[3102] = 8'hdf ;
            rom[3103] = 8'h15 ;
            rom[3104] = 8'h18 ;
            rom[3105] = 8'hf0 ;
            rom[3106] = 8'h07 ;
            rom[3107] = 8'h13 ;
            rom[3108] = 8'h03 ;
            rom[3109] = 8'hfc ;
            rom[3110] = 8'h00 ;
            rom[3111] = 8'hf6 ;
            rom[3112] = 8'h1d ;
            rom[3113] = 8'h0a ;
            rom[3114] = 8'h04 ;
            rom[3115] = 8'h10 ;
            rom[3116] = 8'h39 ;
            rom[3117] = 8'h24 ;
            rom[3118] = 8'h05 ;
            rom[3119] = 8'hee ;
            rom[3120] = 8'hdd ;
            rom[3121] = 8'h4f ;
            rom[3122] = 8'hf2 ;
            rom[3123] = 8'h04 ;
            rom[3124] = 8'h14 ;
            rom[3125] = 8'h24 ;
            rom[3126] = 8'he9 ;
            rom[3127] = 8'hf2 ;
            rom[3128] = 8'hf6 ;
            rom[3129] = 8'hf7 ;
            rom[3130] = 8'h03 ;
            rom[3131] = 8'h03 ;
            rom[3132] = 8'h0b ;
            rom[3133] = 8'hfc ;
            rom[3134] = 8'h0b ;
            rom[3135] = 8'hfd ;
            rom[3136] = 8'h07 ;
            rom[3137] = 8'h11 ;
            rom[3138] = 8'h02 ;
            rom[3139] = 8'hff ;
            rom[3140] = 8'h02 ;
            rom[3141] = 8'hea ;
            rom[3142] = 8'h01 ;
            rom[3143] = 8'h15 ;
            rom[3144] = 8'h1d ;
            rom[3145] = 8'hf0 ;
            rom[3146] = 8'hd5 ;
            rom[3147] = 8'hed ;
            rom[3148] = 8'hf6 ;
            rom[3149] = 8'hfd ;
            rom[3150] = 8'h14 ;
            rom[3151] = 8'h33 ;
            rom[3152] = 8'he5 ;
            rom[3153] = 8'hef ;
            rom[3154] = 8'h07 ;
            rom[3155] = 8'hd4 ;
            rom[3156] = 8'hec ;
            rom[3157] = 8'he6 ;
            rom[3158] = 8'hff ;
            rom[3159] = 8'hdb ;
            rom[3160] = 8'h23 ;
            rom[3161] = 8'h1b ;
            rom[3162] = 8'hfa ;
            rom[3163] = 8'h14 ;
            rom[3164] = 8'h05 ;
            rom[3165] = 8'hf9 ;
            rom[3166] = 8'hf6 ;
            rom[3167] = 8'h19 ;
            rom[3168] = 8'h0e ;
            rom[3169] = 8'h3e ;
            rom[3170] = 8'hf9 ;
            rom[3171] = 8'he7 ;
            rom[3172] = 8'h2c ;
            rom[3173] = 8'hde ;
            rom[3174] = 8'hee ;
            rom[3175] = 8'h25 ;
            rom[3176] = 8'h0f ;
            rom[3177] = 8'h06 ;
            rom[3178] = 8'hf3 ;
            rom[3179] = 8'h20 ;
            rom[3180] = 8'hfa ;
            rom[3181] = 8'hec ;
            rom[3182] = 8'hf9 ;
            rom[3183] = 8'hf1 ;
            rom[3184] = 8'hd9 ;
            rom[3185] = 8'h30 ;
            rom[3186] = 8'h1c ;
            rom[3187] = 8'he4 ;
            rom[3188] = 8'h00 ;
            rom[3189] = 8'hd6 ;
            rom[3190] = 8'h17 ;
            rom[3191] = 8'hfa ;
            rom[3192] = 8'h2e ;
            rom[3193] = 8'h11 ;
            rom[3194] = 8'h0d ;
            rom[3195] = 8'hdb ;
            rom[3196] = 8'hfd ;
            rom[3197] = 8'he2 ;
            rom[3198] = 8'h05 ;
            rom[3199] = 8'hf8 ;
            rom[3200] = 8'hc3 ;
            rom[3201] = 8'h02 ;
            rom[3202] = 8'hfa ;
            rom[3203] = 8'hef ;
            rom[3204] = 8'h01 ;
            rom[3205] = 8'h04 ;
            rom[3206] = 8'hd3 ;
            rom[3207] = 8'hf0 ;
            rom[3208] = 8'h0b ;
            rom[3209] = 8'h14 ;
            rom[3210] = 8'h16 ;
            rom[3211] = 8'he0 ;
            rom[3212] = 8'h00 ;
            rom[3213] = 8'hdc ;
            rom[3214] = 8'h1a ;
            rom[3215] = 8'hfd ;
            rom[3216] = 8'he8 ;
            rom[3217] = 8'hec ;
            rom[3218] = 8'h17 ;
            rom[3219] = 8'h08 ;
            rom[3220] = 8'hf2 ;
            rom[3221] = 8'h15 ;
            rom[3222] = 8'h23 ;
            rom[3223] = 8'h10 ;
            rom[3224] = 8'he8 ;
            rom[3225] = 8'h0f ;
            rom[3226] = 8'hf1 ;
            rom[3227] = 8'hf2 ;
            rom[3228] = 8'he6 ;
            rom[3229] = 8'h08 ;
            rom[3230] = 8'hfa ;
            rom[3231] = 8'hdf ;
            rom[3232] = 8'hf7 ;
            rom[3233] = 8'h0d ;
            rom[3234] = 8'h00 ;
            rom[3235] = 8'hda ;
            rom[3236] = 8'hea ;
            rom[3237] = 8'hea ;
            rom[3238] = 8'hd5 ;
            rom[3239] = 8'h06 ;
            rom[3240] = 8'hf2 ;
            rom[3241] = 8'hf0 ;
            rom[3242] = 8'h11 ;
            rom[3243] = 8'h10 ;
            rom[3244] = 8'h0a ;
            rom[3245] = 8'he4 ;
            rom[3246] = 8'h15 ;
            rom[3247] = 8'h07 ;
            rom[3248] = 8'hfa ;
            rom[3249] = 8'h13 ;
            rom[3250] = 8'hf2 ;
            rom[3251] = 8'h12 ;
            rom[3252] = 8'hef ;
            rom[3253] = 8'h1d ;
            rom[3254] = 8'hf8 ;
            rom[3255] = 8'hd6 ;
            rom[3256] = 8'hff ;
            rom[3257] = 8'hfb ;
            rom[3258] = 8'he7 ;
            rom[3259] = 8'hd9 ;
            rom[3260] = 8'hf0 ;
            rom[3261] = 8'hdf ;
            rom[3262] = 8'h02 ;
            rom[3263] = 8'hfb ;
            rom[3264] = 8'h19 ;
            rom[3265] = 8'hdf ;
            rom[3266] = 8'h1c ;
            rom[3267] = 8'h18 ;
            rom[3268] = 8'hf8 ;
            rom[3269] = 8'hf8 ;
            rom[3270] = 8'hee ;
            rom[3271] = 8'h0f ;
            rom[3272] = 8'hfa ;
            rom[3273] = 8'hee ;
            rom[3274] = 8'hd1 ;
            rom[3275] = 8'h05 ;
            rom[3276] = 8'h05 ;
            rom[3277] = 8'hf6 ;
            rom[3278] = 8'hef ;
            rom[3279] = 8'h03 ;
            rom[3280] = 8'h22 ;
            rom[3281] = 8'hcd ;
            rom[3282] = 8'h0f ;
            rom[3283] = 8'hf3 ;
            rom[3284] = 8'hf6 ;
            rom[3285] = 8'hce ;
            rom[3286] = 8'hee ;
            rom[3287] = 8'hf4 ;
            rom[3288] = 8'hf1 ;
            rom[3289] = 8'hfc ;
            rom[3290] = 8'hf9 ;
            rom[3291] = 8'hef ;
            rom[3292] = 8'h0b ;
            rom[3293] = 8'hdf ;
            rom[3294] = 8'hd5 ;
            rom[3295] = 8'h01 ;
            rom[3296] = 8'h1f ;
            rom[3297] = 8'h23 ;
            rom[3298] = 8'hdd ;
            rom[3299] = 8'hf4 ;
            rom[3300] = 8'h1d ;
            rom[3301] = 8'hfc ;
            rom[3302] = 8'hfb ;
            rom[3303] = 8'h27 ;
            rom[3304] = 8'hf1 ;
            rom[3305] = 8'h21 ;
            rom[3306] = 8'h06 ;
            rom[3307] = 8'h11 ;
            rom[3308] = 8'h22 ;
            rom[3309] = 8'h05 ;
            rom[3310] = 8'he2 ;
            rom[3311] = 8'hdc ;
            rom[3312] = 8'h18 ;
            rom[3313] = 8'hea ;
            rom[3314] = 8'hfa ;
            rom[3315] = 8'he7 ;
            rom[3316] = 8'hfd ;
            rom[3317] = 8'hde ;
            rom[3318] = 8'h04 ;
            rom[3319] = 8'hfb ;
            rom[3320] = 8'h21 ;
            rom[3321] = 8'h0e ;
            rom[3322] = 8'hf4 ;
            rom[3323] = 8'hd7 ;
            rom[3324] = 8'hfb ;
            rom[3325] = 8'he9 ;
            rom[3326] = 8'h03 ;
            rom[3327] = 8'hd9 ;
            rom[3328] = 8'h09 ;
            rom[3329] = 8'hce ;
            rom[3330] = 8'he6 ;
            rom[3331] = 8'h10 ;
            rom[3332] = 8'hf8 ;
            rom[3333] = 8'h06 ;
            rom[3334] = 8'h04 ;
            rom[3335] = 8'h17 ;
            rom[3336] = 8'hd4 ;
            rom[3337] = 8'h06 ;
            rom[3338] = 8'hf2 ;
            rom[3339] = 8'he0 ;
            rom[3340] = 8'hdc ;
            rom[3341] = 8'hfd ;
            rom[3342] = 8'h03 ;
            rom[3343] = 8'h22 ;
            rom[3344] = 8'h03 ;
            rom[3345] = 8'hf7 ;
            rom[3346] = 8'h08 ;
            rom[3347] = 8'h12 ;
            rom[3348] = 8'h01 ;
            rom[3349] = 8'h0a ;
            rom[3350] = 8'hd2 ;
            rom[3351] = 8'h13 ;
            rom[3352] = 8'hf6 ;
            rom[3353] = 8'hcd ;
            rom[3354] = 8'h07 ;
            rom[3355] = 8'hb9 ;
            rom[3356] = 8'h00 ;
            rom[3357] = 8'hfe ;
            rom[3358] = 8'hf6 ;
            rom[3359] = 8'h0e ;
            rom[3360] = 8'h0b ;
            rom[3361] = 8'h09 ;
            rom[3362] = 8'h04 ;
            rom[3363] = 8'hf6 ;
            rom[3364] = 8'h1e ;
            rom[3365] = 8'h09 ;
            rom[3366] = 8'h05 ;
            rom[3367] = 8'hf6 ;
            rom[3368] = 8'hf0 ;
            rom[3369] = 8'h08 ;
            rom[3370] = 8'he6 ;
            rom[3371] = 8'h19 ;
            rom[3372] = 8'h33 ;
            rom[3373] = 8'h1b ;
            rom[3374] = 8'he0 ;
            rom[3375] = 8'heb ;
            rom[3376] = 8'h07 ;
            rom[3377] = 8'hea ;
            rom[3378] = 8'h03 ;
            rom[3379] = 8'hf3 ;
            rom[3380] = 8'hfc ;
            rom[3381] = 8'hf9 ;
            rom[3382] = 8'h00 ;
            rom[3383] = 8'hfc ;
            rom[3384] = 8'hfd ;
            rom[3385] = 8'heb ;
            rom[3386] = 8'h06 ;
            rom[3387] = 8'h08 ;
            rom[3388] = 8'hf0 ;
            rom[3389] = 8'h0b ;
            rom[3390] = 8'h2c ;
            rom[3391] = 8'hf6 ;
            rom[3392] = 8'h21 ;
            rom[3393] = 8'h43 ;
            rom[3394] = 8'h1d ;
            rom[3395] = 8'hd7 ;
            rom[3396] = 8'h13 ;
            rom[3397] = 8'hee ;
            rom[3398] = 8'h0f ;
            rom[3399] = 8'hfc ;
            rom[3400] = 8'he1 ;
            rom[3401] = 8'h0b ;
            rom[3402] = 8'hf1 ;
            rom[3403] = 8'hdc ;
            rom[3404] = 8'hff ;
            rom[3405] = 8'he7 ;
            rom[3406] = 8'h02 ;
            rom[3407] = 8'h10 ;
            rom[3408] = 8'hec ;
            rom[3409] = 8'hf6 ;
            rom[3410] = 8'hf7 ;
            rom[3411] = 8'h0e ;
            rom[3412] = 8'h29 ;
            rom[3413] = 8'h28 ;
            rom[3414] = 8'hee ;
            rom[3415] = 8'he5 ;
            rom[3416] = 8'hfa ;
            rom[3417] = 8'h02 ;
            rom[3418] = 8'hf6 ;
            rom[3419] = 8'h15 ;
            rom[3420] = 8'hdf ;
            rom[3421] = 8'h04 ;
            rom[3422] = 8'hd5 ;
            rom[3423] = 8'h14 ;
            rom[3424] = 8'h0b ;
            rom[3425] = 8'he2 ;
            rom[3426] = 8'h0c ;
            rom[3427] = 8'hec ;
            rom[3428] = 8'hdb ;
            rom[3429] = 8'hf4 ;
            rom[3430] = 8'h17 ;
            rom[3431] = 8'h09 ;
            rom[3432] = 8'heb ;
            rom[3433] = 8'hf4 ;
            rom[3434] = 8'h24 ;
            rom[3435] = 8'h21 ;
            rom[3436] = 8'hf3 ;
            rom[3437] = 8'hc7 ;
            rom[3438] = 8'h08 ;
            rom[3439] = 8'h26 ;
            rom[3440] = 8'hf9 ;
            rom[3441] = 8'h20 ;
            rom[3442] = 8'hf5 ;
            rom[3443] = 8'hf3 ;
            rom[3444] = 8'h28 ;
            rom[3445] = 8'hfe ;
            rom[3446] = 8'h00 ;
            rom[3447] = 8'hf5 ;
            rom[3448] = 8'h18 ;
            rom[3449] = 8'h04 ;
            rom[3450] = 8'he9 ;
            rom[3451] = 8'h21 ;
            rom[3452] = 8'hef ;
            rom[3453] = 8'hf2 ;
            rom[3454] = 8'he7 ;
            rom[3455] = 8'h24 ;
            rom[3456] = 8'hf6 ;
            rom[3457] = 8'he8 ;
            rom[3458] = 8'hca ;
            rom[3459] = 8'h2f ;
            rom[3460] = 8'h1b ;
            rom[3461] = 8'hbf ;
            rom[3462] = 8'hdb ;
            rom[3463] = 8'h1e ;
            rom[3464] = 8'he1 ;
            rom[3465] = 8'hee ;
            rom[3466] = 8'h22 ;
            rom[3467] = 8'hb9 ;
            rom[3468] = 8'hdc ;
            rom[3469] = 8'hdf ;
            rom[3470] = 8'h09 ;
            rom[3471] = 8'hc0 ;
            rom[3472] = 8'hf9 ;
            rom[3473] = 8'hd7 ;
            rom[3474] = 8'hf3 ;
            rom[3475] = 8'hd0 ;
            rom[3476] = 8'hfd ;
            rom[3477] = 8'hd1 ;
            rom[3478] = 8'hf7 ;
            rom[3479] = 8'h04 ;
            rom[3480] = 8'hf0 ;
            rom[3481] = 8'h0a ;
            rom[3482] = 8'hf7 ;
            rom[3483] = 8'hff ;
            rom[3484] = 8'h2d ;
            rom[3485] = 8'h27 ;
            rom[3486] = 8'h09 ;
            rom[3487] = 8'h16 ;
            rom[3488] = 8'h00 ;
            rom[3489] = 8'hfe ;
            rom[3490] = 8'he4 ;
            rom[3491] = 8'h2a ;
            rom[3492] = 8'he9 ;
            rom[3493] = 8'h18 ;
            rom[3494] = 8'he2 ;
            rom[3495] = 8'h16 ;
            rom[3496] = 8'hdd ;
            rom[3497] = 8'h1f ;
            rom[3498] = 8'hf9 ;
            rom[3499] = 8'hfd ;
            rom[3500] = 8'h08 ;
            rom[3501] = 8'he7 ;
            rom[3502] = 8'he7 ;
            rom[3503] = 8'hfb ;
            rom[3504] = 8'h0a ;
            rom[3505] = 8'h25 ;
            rom[3506] = 8'hf2 ;
            rom[3507] = 8'hc5 ;
            rom[3508] = 8'h13 ;
            rom[3509] = 8'hed ;
            rom[3510] = 8'h0e ;
            rom[3511] = 8'h0d ;
            rom[3512] = 8'h17 ;
            rom[3513] = 8'h11 ;
            rom[3514] = 8'h2c ;
            rom[3515] = 8'hde ;
            rom[3516] = 8'hfc ;
            rom[3517] = 8'hf6 ;
            rom[3518] = 8'hfa ;
            rom[3519] = 8'he1 ;
            rom[3520] = 8'h21 ;
            rom[3521] = 8'h03 ;
            rom[3522] = 8'he6 ;
            rom[3523] = 8'heb ;
            rom[3524] = 8'hfb ;
            rom[3525] = 8'hea ;
            rom[3526] = 8'hf3 ;
            rom[3527] = 8'hf2 ;
            rom[3528] = 8'h0f ;
            rom[3529] = 8'hf3 ;
            rom[3530] = 8'hdd ;
            rom[3531] = 8'hf8 ;
            rom[3532] = 8'hf6 ;
            rom[3533] = 8'h19 ;
            rom[3534] = 8'he0 ;
            rom[3535] = 8'h18 ;
            rom[3536] = 8'h36 ;
            rom[3537] = 8'hec ;
            rom[3538] = 8'h04 ;
            rom[3539] = 8'h0c ;
            rom[3540] = 8'hfc ;
            rom[3541] = 8'hf5 ;
            rom[3542] = 8'h16 ;
            rom[3543] = 8'he3 ;
            rom[3544] = 8'h1e ;
            rom[3545] = 8'hfa ;
            rom[3546] = 8'h0c ;
            rom[3547] = 8'h16 ;
            rom[3548] = 8'hc3 ;
            rom[3549] = 8'hf3 ;
            rom[3550] = 8'hb9 ;
            rom[3551] = 8'h05 ;
            rom[3552] = 8'hf5 ;
            rom[3553] = 8'h05 ;
            rom[3554] = 8'h05 ;
            rom[3555] = 8'h19 ;
            rom[3556] = 8'hc8 ;
            rom[3557] = 8'h17 ;
            rom[3558] = 8'h1e ;
            rom[3559] = 8'h00 ;
            rom[3560] = 8'hc6 ;
            rom[3561] = 8'hf0 ;
            rom[3562] = 8'h09 ;
            rom[3563] = 8'h0b ;
            rom[3564] = 8'hea ;
            rom[3565] = 8'h0d ;
            rom[3566] = 8'hb5 ;
            rom[3567] = 8'hfb ;
            rom[3568] = 8'he9 ;
            rom[3569] = 8'h04 ;
            rom[3570] = 8'hea ;
            rom[3571] = 8'h02 ;
            rom[3572] = 8'hef ;
            rom[3573] = 8'h33 ;
            rom[3574] = 8'hfe ;
            rom[3575] = 8'h19 ;
            rom[3576] = 8'hf7 ;
            rom[3577] = 8'hee ;
            rom[3578] = 8'hc7 ;
            rom[3579] = 8'h27 ;
            rom[3580] = 8'hda ;
            rom[3581] = 8'h20 ;
            rom[3582] = 8'h1d ;
            rom[3583] = 8'hf2 ;
            rom[3584] = 8'he6 ;
            rom[3585] = 8'hdd ;
            rom[3586] = 8'h2c ;
            rom[3587] = 8'hdf ;
            rom[3588] = 8'h02 ;
            rom[3589] = 8'h1a ;
            rom[3590] = 8'h14 ;
            rom[3591] = 8'hfc ;
            rom[3592] = 8'hf2 ;
            rom[3593] = 8'he3 ;
            rom[3594] = 8'h0d ;
            rom[3595] = 8'hee ;
            rom[3596] = 8'hef ;
            rom[3597] = 8'hce ;
            rom[3598] = 8'h18 ;
            rom[3599] = 8'hf9 ;
            rom[3600] = 8'hd7 ;
            rom[3601] = 8'h20 ;
            rom[3602] = 8'hdd ;
            rom[3603] = 8'h03 ;
            rom[3604] = 8'h11 ;
            rom[3605] = 8'hcc ;
            rom[3606] = 8'h02 ;
            rom[3607] = 8'hf9 ;
            rom[3608] = 8'he2 ;
            rom[3609] = 8'hef ;
            rom[3610] = 8'hf1 ;
            rom[3611] = 8'h99 ;
            rom[3612] = 8'h01 ;
            rom[3613] = 8'hed ;
            rom[3614] = 8'hfc ;
            rom[3615] = 8'h1b ;
            rom[3616] = 8'h17 ;
            rom[3617] = 8'h1d ;
            rom[3618] = 8'h21 ;
            rom[3619] = 8'hff ;
            rom[3620] = 8'h15 ;
            rom[3621] = 8'hf0 ;
            rom[3622] = 8'h15 ;
            rom[3623] = 8'he0 ;
            rom[3624] = 8'h16 ;
            rom[3625] = 8'hec ;
            rom[3626] = 8'hfb ;
            rom[3627] = 8'h0c ;
            rom[3628] = 8'hee ;
            rom[3629] = 8'hce ;
            rom[3630] = 8'hfc ;
            rom[3631] = 8'h0a ;
            rom[3632] = 8'hbf ;
            rom[3633] = 8'he8 ;
            rom[3634] = 8'hec ;
            rom[3635] = 8'hf6 ;
            rom[3636] = 8'h08 ;
            rom[3637] = 8'hea ;
            rom[3638] = 8'h0b ;
            rom[3639] = 8'h05 ;
            rom[3640] = 8'he8 ;
            rom[3641] = 8'he0 ;
            rom[3642] = 8'h08 ;
            rom[3643] = 8'hf8 ;
            rom[3644] = 8'h11 ;
            rom[3645] = 8'h19 ;
            rom[3646] = 8'h00 ;
            rom[3647] = 8'h10 ;
            rom[3648] = 8'hde ;
            rom[3649] = 8'h12 ;
            rom[3650] = 8'h0c ;
            rom[3651] = 8'h21 ;
            rom[3652] = 8'h08 ;
            rom[3653] = 8'hf7 ;
            rom[3654] = 8'h10 ;
            rom[3655] = 8'h12 ;
            rom[3656] = 8'hf2 ;
            rom[3657] = 8'h07 ;
            rom[3658] = 8'hec ;
            rom[3659] = 8'hfc ;
            rom[3660] = 8'hda ;
            rom[3661] = 8'hd6 ;
            rom[3662] = 8'h03 ;
            rom[3663] = 8'h06 ;
            rom[3664] = 8'hf7 ;
            rom[3665] = 8'hff ;
            rom[3666] = 8'h14 ;
            rom[3667] = 8'hcc ;
            rom[3668] = 8'h03 ;
            rom[3669] = 8'h07 ;
            rom[3670] = 8'he0 ;
            rom[3671] = 8'h30 ;
            rom[3672] = 8'hef ;
            rom[3673] = 8'h06 ;
            rom[3674] = 8'he2 ;
            rom[3675] = 8'h18 ;
            rom[3676] = 8'hc4 ;
            rom[3677] = 8'he9 ;
            rom[3678] = 8'hfd ;
            rom[3679] = 8'h18 ;
            rom[3680] = 8'hcf ;
            rom[3681] = 8'h04 ;
            rom[3682] = 8'hcb ;
            rom[3683] = 8'hf9 ;
            rom[3684] = 8'hf8 ;
            rom[3685] = 8'hfb ;
            rom[3686] = 8'h15 ;
            rom[3687] = 8'h0e ;
            rom[3688] = 8'h11 ;
            rom[3689] = 8'hfb ;
            rom[3690] = 8'h12 ;
            rom[3691] = 8'hf2 ;
            rom[3692] = 8'h07 ;
            rom[3693] = 8'hf1 ;
            rom[3694] = 8'h1b ;
            rom[3695] = 8'hd2 ;
            rom[3696] = 8'hdd ;
            rom[3697] = 8'hf7 ;
            rom[3698] = 8'h10 ;
            rom[3699] = 8'hec ;
            rom[3700] = 8'h0f ;
            rom[3701] = 8'h1e ;
            rom[3702] = 8'hf4 ;
            rom[3703] = 8'h0b ;
            rom[3704] = 8'h14 ;
            rom[3705] = 8'hd6 ;
            rom[3706] = 8'h12 ;
            rom[3707] = 8'hfe ;
            rom[3708] = 8'hf9 ;
            rom[3709] = 8'h1e ;
            rom[3710] = 8'hf9 ;
            rom[3711] = 8'hcc ;
            rom[3712] = 8'hee ;
            rom[3713] = 8'hf5 ;
            rom[3714] = 8'hc5 ;
            rom[3715] = 8'hfc ;
            rom[3716] = 8'hfc ;
            rom[3717] = 8'h0a ;
            rom[3718] = 8'h17 ;
            rom[3719] = 8'h0d ;
            rom[3720] = 8'h12 ;
            rom[3721] = 8'h04 ;
            rom[3722] = 8'he0 ;
            rom[3723] = 8'h08 ;
            rom[3724] = 8'hc9 ;
            rom[3725] = 8'hec ;
            rom[3726] = 8'he5 ;
            rom[3727] = 8'h0a ;
            rom[3728] = 8'h0a ;
            rom[3729] = 8'hee ;
            rom[3730] = 8'h03 ;
            rom[3731] = 8'h0e ;
            rom[3732] = 8'hfe ;
            rom[3733] = 8'h00 ;
            rom[3734] = 8'h07 ;
            rom[3735] = 8'h04 ;
            rom[3736] = 8'hf0 ;
            rom[3737] = 8'h03 ;
            rom[3738] = 8'h06 ;
            rom[3739] = 8'he6 ;
            rom[3740] = 8'h0f ;
            rom[3741] = 8'hfd ;
            rom[3742] = 8'hf0 ;
            rom[3743] = 8'h0f ;
            rom[3744] = 8'h1a ;
            rom[3745] = 8'h20 ;
            rom[3746] = 8'hf3 ;
            rom[3747] = 8'hee ;
            rom[3748] = 8'hd5 ;
            rom[3749] = 8'h16 ;
            rom[3750] = 8'he8 ;
            rom[3751] = 8'h16 ;
            rom[3752] = 8'hd9 ;
            rom[3753] = 8'heb ;
            rom[3754] = 8'hfa ;
            rom[3755] = 8'h10 ;
            rom[3756] = 8'he3 ;
            rom[3757] = 8'h04 ;
            rom[3758] = 8'hef ;
            rom[3759] = 8'h09 ;
            rom[3760] = 8'h05 ;
            rom[3761] = 8'h0d ;
            rom[3762] = 8'he5 ;
            rom[3763] = 8'h06 ;
            rom[3764] = 8'hfa ;
            rom[3765] = 8'hdc ;
            rom[3766] = 8'heb ;
            rom[3767] = 8'hfa ;
            rom[3768] = 8'h0c ;
            rom[3769] = 8'hef ;
            rom[3770] = 8'hf9 ;
            rom[3771] = 8'he3 ;
            rom[3772] = 8'h06 ;
            rom[3773] = 8'hf2 ;
            rom[3774] = 8'hf8 ;
            rom[3775] = 8'he1 ;
            rom[3776] = 8'hea ;
            rom[3777] = 8'hd5 ;
            rom[3778] = 8'h16 ;
            rom[3779] = 8'h07 ;
            rom[3780] = 8'heb ;
            rom[3781] = 8'h0a ;
            rom[3782] = 8'he7 ;
            rom[3783] = 8'he0 ;
            rom[3784] = 8'he0 ;
            rom[3785] = 8'h0f ;
            rom[3786] = 8'hd9 ;
            rom[3787] = 8'hde ;
            rom[3788] = 8'hfe ;
            rom[3789] = 8'h1a ;
            rom[3790] = 8'he8 ;
            rom[3791] = 8'h3d ;
            rom[3792] = 8'h20 ;
            rom[3793] = 8'hfe ;
            rom[3794] = 8'hea ;
            rom[3795] = 8'hfd ;
            rom[3796] = 8'hf5 ;
            rom[3797] = 8'hea ;
            rom[3798] = 8'hf2 ;
            rom[3799] = 8'hc0 ;
            rom[3800] = 8'h04 ;
            rom[3801] = 8'he9 ;
            rom[3802] = 8'hdc ;
            rom[3803] = 8'hf1 ;
            rom[3804] = 8'hf6 ;
            rom[3805] = 8'hef ;
            rom[3806] = 8'hef ;
            rom[3807] = 8'hf2 ;
            rom[3808] = 8'h03 ;
            rom[3809] = 8'hfc ;
            rom[3810] = 8'hcf ;
            rom[3811] = 8'heb ;
            rom[3812] = 8'h04 ;
            rom[3813] = 8'hff ;
            rom[3814] = 8'hfc ;
            rom[3815] = 8'hec ;
            rom[3816] = 8'he9 ;
            rom[3817] = 8'hee ;
            rom[3818] = 8'hfb ;
            rom[3819] = 8'hd7 ;
            rom[3820] = 8'h0d ;
            rom[3821] = 8'hde ;
            rom[3822] = 8'hfd ;
            rom[3823] = 8'he1 ;
            rom[3824] = 8'hf4 ;
            rom[3825] = 8'hef ;
            rom[3826] = 8'h13 ;
            rom[3827] = 8'he6 ;
            rom[3828] = 8'hfc ;
            rom[3829] = 8'hde ;
            rom[3830] = 8'he0 ;
            rom[3831] = 8'hd8 ;
            rom[3832] = 8'hde ;
            rom[3833] = 8'hec ;
            rom[3834] = 8'h11 ;
            rom[3835] = 8'h05 ;
            rom[3836] = 8'hf7 ;
            rom[3837] = 8'he1 ;
            rom[3838] = 8'h20 ;
            rom[3839] = 8'hf1 ;
            rom[3840] = 8'hdb ;
            rom[3841] = 8'h10 ;
            rom[3842] = 8'hfe ;
            rom[3843] = 8'h1f ;
            rom[3844] = 8'hf2 ;
            rom[3845] = 8'hfb ;
            rom[3846] = 8'hf0 ;
            rom[3847] = 8'h1c ;
            rom[3848] = 8'hfe ;
            rom[3849] = 8'h24 ;
            rom[3850] = 8'h00 ;
            rom[3851] = 8'h01 ;
            rom[3852] = 8'hed ;
            rom[3853] = 8'hfa ;
            rom[3854] = 8'he9 ;
            rom[3855] = 8'h0d ;
            rom[3856] = 8'hf9 ;
            rom[3857] = 8'he8 ;
            rom[3858] = 8'h0e ;
            rom[3859] = 8'h05 ;
            rom[3860] = 8'h0c ;
            rom[3861] = 8'h10 ;
            rom[3862] = 8'hf8 ;
            rom[3863] = 8'h16 ;
            rom[3864] = 8'h03 ;
            rom[3865] = 8'hfe ;
            rom[3866] = 8'h18 ;
            rom[3867] = 8'h08 ;
            rom[3868] = 8'h04 ;
            rom[3869] = 8'h22 ;
            rom[3870] = 8'h16 ;
            rom[3871] = 8'hf6 ;
            rom[3872] = 8'h09 ;
            rom[3873] = 8'h03 ;
            rom[3874] = 8'h0c ;
            rom[3875] = 8'h1f ;
            rom[3876] = 8'hec ;
            rom[3877] = 8'h11 ;
            rom[3878] = 8'hcd ;
            rom[3879] = 8'h14 ;
            rom[3880] = 8'hfd ;
            rom[3881] = 8'he9 ;
            rom[3882] = 8'h01 ;
            rom[3883] = 8'hed ;
            rom[3884] = 8'he0 ;
            rom[3885] = 8'he6 ;
            rom[3886] = 8'h1e ;
            rom[3887] = 8'h0a ;
            rom[3888] = 8'h26 ;
            rom[3889] = 8'h11 ;
            rom[3890] = 8'h06 ;
            rom[3891] = 8'he5 ;
            rom[3892] = 8'hda ;
            rom[3893] = 8'hec ;
            rom[3894] = 8'h06 ;
            rom[3895] = 8'h02 ;
            rom[3896] = 8'h26 ;
            rom[3897] = 8'hfc ;
            rom[3898] = 8'h13 ;
            rom[3899] = 8'he4 ;
            rom[3900] = 8'hff ;
            rom[3901] = 8'hee ;
            rom[3902] = 8'hde ;
            rom[3903] = 8'hfb ;
            rom[3904] = 8'h07 ;
            rom[3905] = 8'he6 ;
            rom[3906] = 8'hdc ;
            rom[3907] = 8'hfe ;
            rom[3908] = 8'h0f ;
            rom[3909] = 8'h19 ;
            rom[3910] = 8'he7 ;
            rom[3911] = 8'hf3 ;
            rom[3912] = 8'h1d ;
            rom[3913] = 8'he7 ;
            rom[3914] = 8'hf7 ;
            rom[3915] = 8'h0e ;
            rom[3916] = 8'hef ;
            rom[3917] = 8'h1f ;
            rom[3918] = 8'hc2 ;
            rom[3919] = 8'hbd ;
            rom[3920] = 8'h1a ;
            rom[3921] = 8'hff ;
            rom[3922] = 8'hf6 ;
            rom[3923] = 8'h15 ;
            rom[3924] = 8'hcf ;
            rom[3925] = 8'heb ;
            rom[3926] = 8'hfd ;
            rom[3927] = 8'hd7 ;
            rom[3928] = 8'hf2 ;
            rom[3929] = 8'h05 ;
            rom[3930] = 8'h09 ;
            rom[3931] = 8'hd9 ;
            rom[3932] = 8'hf2 ;
            rom[3933] = 8'hf7 ;
            rom[3934] = 8'hdf ;
            rom[3935] = 8'hd3 ;
            rom[3936] = 8'h04 ;
            rom[3937] = 8'h1d ;
            rom[3938] = 8'hd0 ;
            rom[3939] = 8'h01 ;
            rom[3940] = 8'hf9 ;
            rom[3941] = 8'h17 ;
            rom[3942] = 8'heb ;
            rom[3943] = 8'h0c ;
            rom[3944] = 8'hfd ;
            rom[3945] = 8'hf5 ;
            rom[3946] = 8'hfb ;
            rom[3947] = 8'hd6 ;
            rom[3948] = 8'he1 ;
            rom[3949] = 8'h06 ;
            rom[3950] = 8'hf7 ;
            rom[3951] = 8'hec ;
            rom[3952] = 8'hee ;
            rom[3953] = 8'hf9 ;
            rom[3954] = 8'h02 ;
            rom[3955] = 8'hee ;
            rom[3956] = 8'hf5 ;
            rom[3957] = 8'hff ;
            rom[3958] = 8'h00 ;
            rom[3959] = 8'hf6 ;
            rom[3960] = 8'hdb ;
            rom[3961] = 8'h0d ;
            rom[3962] = 8'hde ;
            rom[3963] = 8'h1b ;
            rom[3964] = 8'he9 ;
            rom[3965] = 8'hf3 ;
            rom[3966] = 8'h2e ;
            rom[3967] = 8'h05 ;
            rom[3968] = 8'hec ;
            rom[3969] = 8'hd0 ;
            rom[3970] = 8'h19 ;
            rom[3971] = 8'hd5 ;
            rom[3972] = 8'hf3 ;
            rom[3973] = 8'h01 ;
            rom[3974] = 8'hf7 ;
            rom[3975] = 8'hfb ;
            rom[3976] = 8'hf6 ;
            rom[3977] = 8'hf7 ;
            rom[3978] = 8'hf0 ;
            rom[3979] = 8'h0b ;
            rom[3980] = 8'h00 ;
            rom[3981] = 8'hef ;
            rom[3982] = 8'hf4 ;
            rom[3983] = 8'h08 ;
            rom[3984] = 8'hea ;
            rom[3985] = 8'hf5 ;
            rom[3986] = 8'hf8 ;
            rom[3987] = 8'hfe ;
            rom[3988] = 8'he6 ;
            rom[3989] = 8'hce ;
            rom[3990] = 8'hd1 ;
            rom[3991] = 8'hf9 ;
            rom[3992] = 8'hca ;
            rom[3993] = 8'hee ;
            rom[3994] = 8'hde ;
            rom[3995] = 8'hca ;
            rom[3996] = 8'h12 ;
            rom[3997] = 8'hdf ;
            rom[3998] = 8'he3 ;
            rom[3999] = 8'hfb ;
            rom[4000] = 8'he0 ;
            rom[4001] = 8'hf1 ;
            rom[4002] = 8'hee ;
            rom[4003] = 8'hf8 ;
            rom[4004] = 8'he9 ;
            rom[4005] = 8'hf2 ;
            rom[4006] = 8'hf2 ;
            rom[4007] = 8'h11 ;
            rom[4008] = 8'h05 ;
            rom[4009] = 8'hed ;
            rom[4010] = 8'h29 ;
            rom[4011] = 8'hdd ;
            rom[4012] = 8'hc3 ;
            rom[4013] = 8'hc9 ;
            rom[4014] = 8'hee ;
            rom[4015] = 8'hed ;
            rom[4016] = 8'h1b ;
            rom[4017] = 8'hea ;
            rom[4018] = 8'hee ;
            rom[4019] = 8'he5 ;
            rom[4020] = 8'h10 ;
            rom[4021] = 8'h0a ;
            rom[4022] = 8'hfa ;
            rom[4023] = 8'h02 ;
            rom[4024] = 8'he8 ;
            rom[4025] = 8'h0e ;
            rom[4026] = 8'hc6 ;
            rom[4027] = 8'hed ;
            rom[4028] = 8'hfa ;
            rom[4029] = 8'hf5 ;
            rom[4030] = 8'h11 ;
            rom[4031] = 8'hd0 ;
            rom[4032] = 8'hea ;
            rom[4033] = 8'hfb ;
            rom[4034] = 8'hf1 ;
            rom[4035] = 8'hf9 ;
            rom[4036] = 8'h07 ;
            rom[4037] = 8'hf1 ;
            rom[4038] = 8'he7 ;
            rom[4039] = 8'hf3 ;
            rom[4040] = 8'hda ;
            rom[4041] = 8'hee ;
            rom[4042] = 8'h05 ;
            rom[4043] = 8'h08 ;
            rom[4044] = 8'hf1 ;
            rom[4045] = 8'hf3 ;
            rom[4046] = 8'h17 ;
            rom[4047] = 8'he7 ;
            rom[4048] = 8'h01 ;
            rom[4049] = 8'h04 ;
            rom[4050] = 8'he6 ;
            rom[4051] = 8'hff ;
            rom[4052] = 8'h0f ;
            rom[4053] = 8'he3 ;
            rom[4054] = 8'hee ;
            rom[4055] = 8'h15 ;
            rom[4056] = 8'hea ;
            rom[4057] = 8'he2 ;
            rom[4058] = 8'hfb ;
            rom[4059] = 8'h16 ;
            rom[4060] = 8'hdb ;
            rom[4061] = 8'hcf ;
            rom[4062] = 8'h02 ;
            rom[4063] = 8'hff ;
            rom[4064] = 8'hcb ;
            rom[4065] = 8'hdf ;
            rom[4066] = 8'hff ;
            rom[4067] = 8'h0e ;
            rom[4068] = 8'hec ;
            rom[4069] = 8'h0a ;
            rom[4070] = 8'he6 ;
            rom[4071] = 8'hde ;
            rom[4072] = 8'he1 ;
            rom[4073] = 8'hfd ;
            rom[4074] = 8'he9 ;
            rom[4075] = 8'h1d ;
            rom[4076] = 8'h0b ;
            rom[4077] = 8'hfb ;
            rom[4078] = 8'h16 ;
            rom[4079] = 8'hfd ;
            rom[4080] = 8'hd6 ;
            rom[4081] = 8'hfa ;
            rom[4082] = 8'h10 ;
            rom[4083] = 8'hff ;
            rom[4084] = 8'hdd ;
            rom[4085] = 8'h1e ;
            rom[4086] = 8'he0 ;
            rom[4087] = 8'hfb ;
            rom[4088] = 8'hf4 ;
            rom[4089] = 8'hd5 ;
            rom[4090] = 8'hed ;
            rom[4091] = 8'he7 ;
            rom[4092] = 8'h08 ;
            rom[4093] = 8'hf4 ;
            rom[4094] = 8'he6 ;
            rom[4095] = 8'hf6 ;
            rom[4096] = 8'h01 ;
            rom[4097] = 8'h19 ;
            rom[4098] = 8'hc6 ;
            rom[4099] = 8'h1f ;
            rom[4100] = 8'h1e ;
            rom[4101] = 8'h08 ;
            rom[4102] = 8'hec ;
            rom[4103] = 8'heb ;
            rom[4104] = 8'h15 ;
            rom[4105] = 8'hfa ;
            rom[4106] = 8'hf5 ;
            rom[4107] = 8'he9 ;
            rom[4108] = 8'hf0 ;
            rom[4109] = 8'hfc ;
            rom[4110] = 8'h07 ;
            rom[4111] = 8'hb6 ;
            rom[4112] = 8'h19 ;
            rom[4113] = 8'he2 ;
            rom[4114] = 8'h01 ;
            rom[4115] = 8'h03 ;
            rom[4116] = 8'h0a ;
            rom[4117] = 8'hf5 ;
            rom[4118] = 8'h13 ;
            rom[4119] = 8'h1a ;
            rom[4120] = 8'hf6 ;
            rom[4121] = 8'h14 ;
            rom[4122] = 8'h0b ;
            rom[4123] = 8'heb ;
            rom[4124] = 8'h1a ;
            rom[4125] = 8'h1a ;
            rom[4126] = 8'hf8 ;
            rom[4127] = 8'h1a ;
            rom[4128] = 8'h10 ;
            rom[4129] = 8'h1d ;
            rom[4130] = 8'h06 ;
            rom[4131] = 8'hfa ;
            rom[4132] = 8'he6 ;
            rom[4133] = 8'hd5 ;
            rom[4134] = 8'hbc ;
            rom[4135] = 8'h1e ;
            rom[4136] = 8'hea ;
            rom[4137] = 8'he2 ;
            rom[4138] = 8'hdd ;
            rom[4139] = 8'h09 ;
            rom[4140] = 8'h00 ;
            rom[4141] = 8'hec ;
            rom[4142] = 8'hf9 ;
            rom[4143] = 8'he0 ;
            rom[4144] = 8'h19 ;
            rom[4145] = 8'h1f ;
            rom[4146] = 8'hcf ;
            rom[4147] = 8'he8 ;
            rom[4148] = 8'hc4 ;
            rom[4149] = 8'hf8 ;
            rom[4150] = 8'h0a ;
            rom[4151] = 8'h0c ;
            rom[4152] = 8'h0a ;
            rom[4153] = 8'hf0 ;
            rom[4154] = 8'h1d ;
            rom[4155] = 8'hdc ;
            rom[4156] = 8'hed ;
            rom[4157] = 8'hdb ;
            rom[4158] = 8'he9 ;
            rom[4159] = 8'hf2 ;
            rom[4160] = 8'h05 ;
            rom[4161] = 8'he3 ;
            rom[4162] = 8'h17 ;
            rom[4163] = 8'hf5 ;
            rom[4164] = 8'h11 ;
            rom[4165] = 8'h25 ;
            rom[4166] = 8'hfa ;
            rom[4167] = 8'hdf ;
            rom[4168] = 8'h0a ;
            rom[4169] = 8'hdc ;
            rom[4170] = 8'he0 ;
            rom[4171] = 8'heb ;
            rom[4172] = 8'hf7 ;
            rom[4173] = 8'hda ;
            rom[4174] = 8'hc9 ;
            rom[4175] = 8'h03 ;
            rom[4176] = 8'h2e ;
            rom[4177] = 8'hc4 ;
            rom[4178] = 8'h0d ;
            rom[4179] = 8'hf8 ;
            rom[4180] = 8'hec ;
            rom[4181] = 8'h13 ;
            rom[4182] = 8'hde ;
            rom[4183] = 8'he9 ;
            rom[4184] = 8'he3 ;
            rom[4185] = 8'h1b ;
            rom[4186] = 8'h19 ;
            rom[4187] = 8'hfb ;
            rom[4188] = 8'hdd ;
            rom[4189] = 8'h05 ;
            rom[4190] = 8'h08 ;
            rom[4191] = 8'hcc ;
            rom[4192] = 8'h17 ;
            rom[4193] = 8'hf4 ;
            rom[4194] = 8'h00 ;
            rom[4195] = 8'h23 ;
            rom[4196] = 8'he7 ;
            rom[4197] = 8'h15 ;
            rom[4198] = 8'h25 ;
            rom[4199] = 8'h0d ;
            rom[4200] = 8'hf3 ;
            rom[4201] = 8'heb ;
            rom[4202] = 8'h1d ;
            rom[4203] = 8'hef ;
            rom[4204] = 8'h0d ;
            rom[4205] = 8'h18 ;
            rom[4206] = 8'hdb ;
            rom[4207] = 8'he9 ;
            rom[4208] = 8'hf8 ;
            rom[4209] = 8'hed ;
            rom[4210] = 8'h06 ;
            rom[4211] = 8'he4 ;
            rom[4212] = 8'hf2 ;
            rom[4213] = 8'hdf ;
            rom[4214] = 8'hd7 ;
            rom[4215] = 8'hef ;
            rom[4216] = 8'hcd ;
            rom[4217] = 8'hf1 ;
            rom[4218] = 8'he5 ;
            rom[4219] = 8'h2c ;
            rom[4220] = 8'hd0 ;
            rom[4221] = 8'h0d ;
            rom[4222] = 8'h09 ;
            rom[4223] = 8'hf6 ;
            rom[4224] = 8'hed ;
            rom[4225] = 8'hd1 ;
            rom[4226] = 8'h20 ;
            rom[4227] = 8'he8 ;
            rom[4228] = 8'h0c ;
            rom[4229] = 8'hfc ;
            rom[4230] = 8'hd0 ;
            rom[4231] = 8'hf7 ;
            rom[4232] = 8'hf0 ;
            rom[4233] = 8'h00 ;
            rom[4234] = 8'h0c ;
            rom[4235] = 8'hf1 ;
            rom[4236] = 8'hf4 ;
            rom[4237] = 8'h03 ;
            rom[4238] = 8'h00 ;
            rom[4239] = 8'h07 ;
            rom[4240] = 8'hed ;
            rom[4241] = 8'h22 ;
            rom[4242] = 8'hee ;
            rom[4243] = 8'hfc ;
            rom[4244] = 8'h07 ;
            rom[4245] = 8'hce ;
            rom[4246] = 8'h13 ;
            rom[4247] = 8'h11 ;
            rom[4248] = 8'he6 ;
            rom[4249] = 8'hf5 ;
            rom[4250] = 8'h17 ;
            rom[4251] = 8'he0 ;
            rom[4252] = 8'hef ;
            rom[4253] = 8'h0f ;
            rom[4254] = 8'h24 ;
            rom[4255] = 8'h18 ;
            rom[4256] = 8'h04 ;
            rom[4257] = 8'h02 ;
            rom[4258] = 8'hcc ;
            rom[4259] = 8'he5 ;
            rom[4260] = 8'hfc ;
            rom[4261] = 8'hf5 ;
            rom[4262] = 8'h17 ;
            rom[4263] = 8'h03 ;
            rom[4264] = 8'hfa ;
            rom[4265] = 8'he9 ;
            rom[4266] = 8'hd2 ;
            rom[4267] = 8'hf4 ;
            rom[4268] = 8'h03 ;
            rom[4269] = 8'he8 ;
            rom[4270] = 8'hf9 ;
            rom[4271] = 8'he5 ;
            rom[4272] = 8'hec ;
            rom[4273] = 8'hca ;
            rom[4274] = 8'hf2 ;
            rom[4275] = 8'hc8 ;
            rom[4276] = 8'h07 ;
            rom[4277] = 8'hf1 ;
            rom[4278] = 8'h1e ;
            rom[4279] = 8'hfa ;
            rom[4280] = 8'h0a ;
            rom[4281] = 8'h0d ;
            rom[4282] = 8'hf8 ;
            rom[4283] = 8'hd7 ;
            rom[4284] = 8'h31 ;
            rom[4285] = 8'h01 ;
            rom[4286] = 8'h27 ;
            rom[4287] = 8'hf7 ;
            rom[4288] = 8'hf6 ;
            rom[4289] = 8'hf2 ;
            rom[4290] = 8'h26 ;
            rom[4291] = 8'h02 ;
            rom[4292] = 8'he5 ;
            rom[4293] = 8'hdd ;
            rom[4294] = 8'h0d ;
            rom[4295] = 8'he2 ;
            rom[4296] = 8'hd7 ;
            rom[4297] = 8'h0b ;
            rom[4298] = 8'h19 ;
            rom[4299] = 8'h14 ;
            rom[4300] = 8'hfe ;
            rom[4301] = 8'hff ;
            rom[4302] = 8'hd8 ;
            rom[4303] = 8'h28 ;
            rom[4304] = 8'hd5 ;
            rom[4305] = 8'hf4 ;
            rom[4306] = 8'h02 ;
            rom[4307] = 8'hf9 ;
            rom[4308] = 8'h02 ;
            rom[4309] = 8'hf4 ;
            rom[4310] = 8'h0f ;
            rom[4311] = 8'h1c ;
            rom[4312] = 8'hef ;
            rom[4313] = 8'hf5 ;
            rom[4314] = 8'hd6 ;
            rom[4315] = 8'h1b ;
            rom[4316] = 8'h01 ;
            rom[4317] = 8'h08 ;
            rom[4318] = 8'h08 ;
            rom[4319] = 8'hf0 ;
            rom[4320] = 8'h08 ;
            rom[4321] = 8'hf3 ;
            rom[4322] = 8'h1d ;
            rom[4323] = 8'hf3 ;
            rom[4324] = 8'hcc ;
            rom[4325] = 8'hd9 ;
            rom[4326] = 8'h0c ;
            rom[4327] = 8'hfb ;
            rom[4328] = 8'hfb ;
            rom[4329] = 8'h11 ;
            rom[4330] = 8'hdc ;
            rom[4331] = 8'hff ;
            rom[4332] = 8'h1e ;
            rom[4333] = 8'h10 ;
            rom[4334] = 8'h0a ;
            rom[4335] = 8'h22 ;
            rom[4336] = 8'h00 ;
            rom[4337] = 8'hf4 ;
            rom[4338] = 8'hf8 ;
            rom[4339] = 8'h11 ;
            rom[4340] = 8'h09 ;
            rom[4341] = 8'hb4 ;
            rom[4342] = 8'h19 ;
            rom[4343] = 8'h14 ;
            rom[4344] = 8'h10 ;
            rom[4345] = 8'h0c ;
            rom[4346] = 8'h01 ;
            rom[4347] = 8'hd7 ;
            rom[4348] = 8'h09 ;
            rom[4349] = 8'h1a ;
            rom[4350] = 8'hc2 ;
            rom[4351] = 8'h04 ;
            rom[4352] = 8'h0e ;
            rom[4353] = 8'h0f ;
            rom[4354] = 8'hf5 ;
            rom[4355] = 8'h10 ;
            rom[4356] = 8'h0a ;
            rom[4357] = 8'hfe ;
            rom[4358] = 8'hfa ;
            rom[4359] = 8'hd8 ;
            rom[4360] = 8'he9 ;
            rom[4361] = 8'h02 ;
            rom[4362] = 8'h0c ;
            rom[4363] = 8'h15 ;
            rom[4364] = 8'h15 ;
            rom[4365] = 8'hfa ;
            rom[4366] = 8'h0a ;
            rom[4367] = 8'hd7 ;
            rom[4368] = 8'hfa ;
            rom[4369] = 8'hfa ;
            rom[4370] = 8'hfe ;
            rom[4371] = 8'he8 ;
            rom[4372] = 8'hfd ;
            rom[4373] = 8'hf4 ;
            rom[4374] = 8'hf9 ;
            rom[4375] = 8'hff ;
            rom[4376] = 8'h09 ;
            rom[4377] = 8'hf8 ;
            rom[4378] = 8'hfb ;
            rom[4379] = 8'he5 ;
            rom[4380] = 8'hfc ;
            rom[4381] = 8'h24 ;
            rom[4382] = 8'h01 ;
            rom[4383] = 8'h10 ;
            rom[4384] = 8'he8 ;
            rom[4385] = 8'h2b ;
            rom[4386] = 8'h1c ;
            rom[4387] = 8'h19 ;
            rom[4388] = 8'h0b ;
            rom[4389] = 8'h13 ;
            rom[4390] = 8'he8 ;
            rom[4391] = 8'h0b ;
            rom[4392] = 8'hff ;
            rom[4393] = 8'hfa ;
            rom[4394] = 8'hf8 ;
            rom[4395] = 8'h06 ;
            rom[4396] = 8'h27 ;
            rom[4397] = 8'h0b ;
            rom[4398] = 8'h14 ;
            rom[4399] = 8'hcc ;
            rom[4400] = 8'he3 ;
            rom[4401] = 8'h1b ;
            rom[4402] = 8'hc5 ;
            rom[4403] = 8'hd5 ;
            rom[4404] = 8'h0e ;
            rom[4405] = 8'h0e ;
            rom[4406] = 8'he0 ;
            rom[4407] = 8'hfd ;
            rom[4408] = 8'h2d ;
            rom[4409] = 8'hd8 ;
            rom[4410] = 8'hf2 ;
            rom[4411] = 8'h03 ;
            rom[4412] = 8'h29 ;
            rom[4413] = 8'hdc ;
            rom[4414] = 8'h18 ;
            rom[4415] = 8'hec ;
            rom[4416] = 8'h26 ;
            rom[4417] = 8'h04 ;
            rom[4418] = 8'h01 ;
            rom[4419] = 8'h1b ;
            rom[4420] = 8'hf5 ;
            rom[4421] = 8'hfd ;
            rom[4422] = 8'he2 ;
            rom[4423] = 8'hcd ;
            rom[4424] = 8'h06 ;
            rom[4425] = 8'h00 ;
            rom[4426] = 8'hde ;
            rom[4427] = 8'hf1 ;
            rom[4428] = 8'he5 ;
            rom[4429] = 8'h1f ;
            rom[4430] = 8'hfd ;
            rom[4431] = 8'h16 ;
            rom[4432] = 8'hee ;
            rom[4433] = 8'he9 ;
            rom[4434] = 8'h0a ;
            rom[4435] = 8'h16 ;
            rom[4436] = 8'hf6 ;
            rom[4437] = 8'hf1 ;
            rom[4438] = 8'he1 ;
            rom[4439] = 8'hde ;
            rom[4440] = 8'hf3 ;
            rom[4441] = 8'h13 ;
            rom[4442] = 8'he8 ;
            rom[4443] = 8'h0c ;
            rom[4444] = 8'hc7 ;
            rom[4445] = 8'h10 ;
            rom[4446] = 8'h09 ;
            rom[4447] = 8'h16 ;
            rom[4448] = 8'h0e ;
            rom[4449] = 8'hff ;
            rom[4450] = 8'hf8 ;
            rom[4451] = 8'h0e ;
            rom[4452] = 8'heb ;
            rom[4453] = 8'hf9 ;
            rom[4454] = 8'heb ;
            rom[4455] = 8'h0a ;
            rom[4456] = 8'hf6 ;
            rom[4457] = 8'hda ;
            rom[4458] = 8'h09 ;
            rom[4459] = 8'h0a ;
            rom[4460] = 8'h00 ;
            rom[4461] = 8'hde ;
            rom[4462] = 8'h15 ;
            rom[4463] = 8'hee ;
            rom[4464] = 8'hca ;
            rom[4465] = 8'heb ;
            rom[4466] = 8'he2 ;
            rom[4467] = 8'h05 ;
            rom[4468] = 8'h16 ;
            rom[4469] = 8'h18 ;
            rom[4470] = 8'hf8 ;
            rom[4471] = 8'hfb ;
            rom[4472] = 8'heb ;
            rom[4473] = 8'h00 ;
            rom[4474] = 8'h02 ;
            rom[4475] = 8'h20 ;
            rom[4476] = 8'h0b ;
            rom[4477] = 8'h13 ;
            rom[4478] = 8'h07 ;
            rom[4479] = 8'hda ;
            rom[4480] = 8'h11 ;
            rom[4481] = 8'hd0 ;
            rom[4482] = 8'h23 ;
            rom[4483] = 8'hfa ;
            rom[4484] = 8'hfd ;
            rom[4485] = 8'h0c ;
            rom[4486] = 8'h00 ;
            rom[4487] = 8'hdf ;
            rom[4488] = 8'h07 ;
            rom[4489] = 8'hd3 ;
            rom[4490] = 8'he4 ;
            rom[4491] = 8'h16 ;
            rom[4492] = 8'h24 ;
            rom[4493] = 8'he8 ;
            rom[4494] = 8'h01 ;
            rom[4495] = 8'h02 ;
            rom[4496] = 8'he4 ;
            rom[4497] = 8'h20 ;
            rom[4498] = 8'h01 ;
            rom[4499] = 8'h0d ;
            rom[4500] = 8'hed ;
            rom[4501] = 8'hd1 ;
            rom[4502] = 8'h1c ;
            rom[4503] = 8'h14 ;
            rom[4504] = 8'h24 ;
            rom[4505] = 8'hce ;
            rom[4506] = 8'h11 ;
            rom[4507] = 8'hcb ;
            rom[4508] = 8'hdf ;
            rom[4509] = 8'h0e ;
            rom[4510] = 8'h03 ;
            rom[4511] = 8'h0b ;
            rom[4512] = 8'hf7 ;
            rom[4513] = 8'h03 ;
            rom[4514] = 8'he1 ;
            rom[4515] = 8'hfc ;
            rom[4516] = 8'h07 ;
            rom[4517] = 8'h0f ;
            rom[4518] = 8'h00 ;
            rom[4519] = 8'hce ;
            rom[4520] = 8'he1 ;
            rom[4521] = 8'heb ;
            rom[4522] = 8'h07 ;
            rom[4523] = 8'h0d ;
            rom[4524] = 8'h15 ;
            rom[4525] = 8'hed ;
            rom[4526] = 8'hf5 ;
            rom[4527] = 8'h08 ;
            rom[4528] = 8'hcc ;
            rom[4529] = 8'hdb ;
            rom[4530] = 8'he6 ;
            rom[4531] = 8'hf4 ;
            rom[4532] = 8'h04 ;
            rom[4533] = 8'hf2 ;
            rom[4534] = 8'hd5 ;
            rom[4535] = 8'h00 ;
            rom[4536] = 8'h11 ;
            rom[4537] = 8'h0a ;
            rom[4538] = 8'hea ;
            rom[4539] = 8'hf2 ;
            rom[4540] = 8'h31 ;
            rom[4541] = 8'hf9 ;
            rom[4542] = 8'h01 ;
            rom[4543] = 8'hf4 ;
            rom[4544] = 8'he2 ;
            rom[4545] = 8'hfb ;
            rom[4546] = 8'h1a ;
            rom[4547] = 8'h0c ;
            rom[4548] = 8'hf8 ;
            rom[4549] = 8'h03 ;
            rom[4550] = 8'hec ;
            rom[4551] = 8'h00 ;
            rom[4552] = 8'hd6 ;
            rom[4553] = 8'h11 ;
            rom[4554] = 8'he4 ;
            rom[4555] = 8'hd3 ;
            rom[4556] = 8'hdc ;
            rom[4557] = 8'hee ;
            rom[4558] = 8'hf8 ;
            rom[4559] = 8'h08 ;
            rom[4560] = 8'hef ;
            rom[4561] = 8'h18 ;
            rom[4562] = 8'h00 ;
            rom[4563] = 8'hd2 ;
            rom[4564] = 8'hdd ;
            rom[4565] = 8'h0b ;
            rom[4566] = 8'he4 ;
            rom[4567] = 8'h09 ;
            rom[4568] = 8'hfa ;
            rom[4569] = 8'h05 ;
            rom[4570] = 8'hd7 ;
            rom[4571] = 8'heb ;
            rom[4572] = 8'h09 ;
            rom[4573] = 8'hf9 ;
            rom[4574] = 8'h33 ;
            rom[4575] = 8'he7 ;
            rom[4576] = 8'he1 ;
            rom[4577] = 8'h1c ;
            rom[4578] = 8'h0f ;
            rom[4579] = 8'h05 ;
            rom[4580] = 8'hd4 ;
            rom[4581] = 8'hed ;
            rom[4582] = 8'hdd ;
            rom[4583] = 8'h0b ;
            rom[4584] = 8'h16 ;
            rom[4585] = 8'h24 ;
            rom[4586] = 8'hef ;
            rom[4587] = 8'h07 ;
            rom[4588] = 8'h22 ;
            rom[4589] = 8'h00 ;
            rom[4590] = 8'he3 ;
            rom[4591] = 8'hf2 ;
            rom[4592] = 8'he1 ;
            rom[4593] = 8'hfb ;
            rom[4594] = 8'he7 ;
            rom[4595] = 8'hfc ;
            rom[4596] = 8'hf8 ;
            rom[4597] = 8'hea ;
            rom[4598] = 8'hfd ;
            rom[4599] = 8'he7 ;
            rom[4600] = 8'h06 ;
            rom[4601] = 8'hff ;
            rom[4602] = 8'hfd ;
            rom[4603] = 8'hed ;
            rom[4604] = 8'h00 ;
            rom[4605] = 8'h0a ;
            rom[4606] = 8'he9 ;
            rom[4607] = 8'h2e ;
            rom[4608] = 8'h00 ;
            rom[4609] = 8'h12 ;
            rom[4610] = 8'h0b ;
            rom[4611] = 8'hf8 ;
            rom[4612] = 8'h1a ;
            rom[4613] = 8'hf1 ;
            rom[4614] = 8'hf9 ;
            rom[4615] = 8'hf7 ;
            rom[4616] = 8'hee ;
            rom[4617] = 8'h0a ;
            rom[4618] = 8'he0 ;
            rom[4619] = 8'hf9 ;
            rom[4620] = 8'h15 ;
            rom[4621] = 8'h10 ;
            rom[4622] = 8'h00 ;
            rom[4623] = 8'hfe ;
            rom[4624] = 8'he0 ;
            rom[4625] = 8'h18 ;
            rom[4626] = 8'he2 ;
            rom[4627] = 8'hea ;
            rom[4628] = 8'hf4 ;
            rom[4629] = 8'hf7 ;
            rom[4630] = 8'hf1 ;
            rom[4631] = 8'h0e ;
            rom[4632] = 8'h22 ;
            rom[4633] = 8'hf4 ;
            rom[4634] = 8'hf3 ;
            rom[4635] = 8'h02 ;
            rom[4636] = 8'h07 ;
            rom[4637] = 8'hf6 ;
            rom[4638] = 8'hfd ;
            rom[4639] = 8'h0f ;
            rom[4640] = 8'h1d ;
            rom[4641] = 8'hf6 ;
            rom[4642] = 8'he8 ;
            rom[4643] = 8'hee ;
            rom[4644] = 8'hfa ;
            rom[4645] = 8'hed ;
            rom[4646] = 8'hf8 ;
            rom[4647] = 8'hec ;
            rom[4648] = 8'h26 ;
            rom[4649] = 8'hd7 ;
            rom[4650] = 8'hfd ;
            rom[4651] = 8'he1 ;
            rom[4652] = 8'h14 ;
            rom[4653] = 8'hfc ;
            rom[4654] = 8'hc4 ;
            rom[4655] = 8'h04 ;
            rom[4656] = 8'h0d ;
            rom[4657] = 8'hf7 ;
            rom[4658] = 8'h13 ;
            rom[4659] = 8'h0a ;
            rom[4660] = 8'hf8 ;
            rom[4661] = 8'h1d ;
            rom[4662] = 8'he5 ;
            rom[4663] = 8'hd1 ;
            rom[4664] = 8'h07 ;
            rom[4665] = 8'hfc ;
            rom[4666] = 8'hcd ;
            rom[4667] = 8'h1e ;
            rom[4668] = 8'he3 ;
            rom[4669] = 8'hf5 ;
            rom[4670] = 8'hda ;
            rom[4671] = 8'h0b ;
            rom[4672] = 8'hf8 ;
            rom[4673] = 8'hef ;
            rom[4674] = 8'hdd ;
            rom[4675] = 8'hd5 ;
            rom[4676] = 8'hea ;
            rom[4677] = 8'hef ;
            rom[4678] = 8'hdf ;
            rom[4679] = 8'hd2 ;
            rom[4680] = 8'hf8 ;
            rom[4681] = 8'h09 ;
            rom[4682] = 8'hff ;
            rom[4683] = 8'h2a ;
            rom[4684] = 8'hfb ;
            rom[4685] = 8'hec ;
            rom[4686] = 8'hf4 ;
            rom[4687] = 8'hea ;
            rom[4688] = 8'hf1 ;
            rom[4689] = 8'h1c ;
            rom[4690] = 8'hc1 ;
            rom[4691] = 8'hef ;
            rom[4692] = 8'hfb ;
            rom[4693] = 8'hf6 ;
            rom[4694] = 8'h06 ;
            rom[4695] = 8'hea ;
            rom[4696] = 8'hee ;
            rom[4697] = 8'h0a ;
            rom[4698] = 8'hfd ;
            rom[4699] = 8'hfb ;
            rom[4700] = 8'hff ;
            rom[4701] = 8'h10 ;
            rom[4702] = 8'h15 ;
            rom[4703] = 8'he4 ;
            rom[4704] = 8'hff ;
            rom[4705] = 8'h16 ;
            rom[4706] = 8'he9 ;
            rom[4707] = 8'h06 ;
            rom[4708] = 8'h0f ;
            rom[4709] = 8'hf6 ;
            rom[4710] = 8'h12 ;
            rom[4711] = 8'hf9 ;
            rom[4712] = 8'heb ;
            rom[4713] = 8'h09 ;
            rom[4714] = 8'hea ;
            rom[4715] = 8'h10 ;
            rom[4716] = 8'hd6 ;
            rom[4717] = 8'h01 ;
            rom[4718] = 8'he7 ;
            rom[4719] = 8'h1c ;
            rom[4720] = 8'h10 ;
            rom[4721] = 8'h11 ;
            rom[4722] = 8'hfa ;
            rom[4723] = 8'he2 ;
            rom[4724] = 8'hef ;
            rom[4725] = 8'h01 ;
            rom[4726] = 8'h06 ;
            rom[4727] = 8'hfe ;
            rom[4728] = 8'hdb ;
            rom[4729] = 8'hf9 ;
            rom[4730] = 8'hfa ;
            rom[4731] = 8'hf1 ;
            rom[4732] = 8'hd9 ;
            rom[4733] = 8'hc0 ;
            rom[4734] = 8'hc9 ;
            rom[4735] = 8'h05 ;
            rom[4736] = 8'he4 ;
            rom[4737] = 8'h00 ;
            rom[4738] = 8'hfc ;
            rom[4739] = 8'h0f ;
            rom[4740] = 8'h1a ;
            rom[4741] = 8'hf1 ;
            rom[4742] = 8'hfc ;
            rom[4743] = 8'h04 ;
            rom[4744] = 8'heb ;
            rom[4745] = 8'h0d ;
            rom[4746] = 8'h03 ;
            rom[4747] = 8'hea ;
            rom[4748] = 8'h00 ;
            rom[4749] = 8'h14 ;
            rom[4750] = 8'hfd ;
            rom[4751] = 8'hfc ;
            rom[4752] = 8'h04 ;
            rom[4753] = 8'he5 ;
            rom[4754] = 8'hd7 ;
            rom[4755] = 8'he8 ;
            rom[4756] = 8'hf3 ;
            rom[4757] = 8'hed ;
            rom[4758] = 8'h21 ;
            rom[4759] = 8'h0f ;
            rom[4760] = 8'h14 ;
            rom[4761] = 8'hee ;
            rom[4762] = 8'h25 ;
            rom[4763] = 8'h23 ;
            rom[4764] = 8'hf5 ;
            rom[4765] = 8'h03 ;
            rom[4766] = 8'h04 ;
            rom[4767] = 8'hb7 ;
            rom[4768] = 8'h2b ;
            rom[4769] = 8'h07 ;
            rom[4770] = 8'h0f ;
            rom[4771] = 8'hd0 ;
            rom[4772] = 8'h07 ;
            rom[4773] = 8'h1e ;
            rom[4774] = 8'h25 ;
            rom[4775] = 8'h0f ;
            rom[4776] = 8'h18 ;
            rom[4777] = 8'he9 ;
            rom[4778] = 8'hf3 ;
            rom[4779] = 8'h07 ;
            rom[4780] = 8'h04 ;
            rom[4781] = 8'h02 ;
            rom[4782] = 8'h39 ;
            rom[4783] = 8'he9 ;
            rom[4784] = 8'he2 ;
            rom[4785] = 8'h13 ;
            rom[4786] = 8'h0c ;
            rom[4787] = 8'he2 ;
            rom[4788] = 8'hfc ;
            rom[4789] = 8'h04 ;
            rom[4790] = 8'h10 ;
            rom[4791] = 8'hf3 ;
            rom[4792] = 8'h38 ;
            rom[4793] = 8'hd5 ;
            rom[4794] = 8'heb ;
            rom[4795] = 8'h04 ;
            rom[4796] = 8'hd5 ;
            rom[4797] = 8'hf6 ;
            rom[4798] = 8'hcb ;
            rom[4799] = 8'h02 ;
            rom[4800] = 8'h16 ;
            rom[4801] = 8'he5 ;
            rom[4802] = 8'hde ;
            rom[4803] = 8'hf5 ;
            rom[4804] = 8'hfc ;
            rom[4805] = 8'hc2 ;
            rom[4806] = 8'hfb ;
            rom[4807] = 8'hfa ;
            rom[4808] = 8'hf7 ;
            rom[4809] = 8'hef ;
            rom[4810] = 8'h0d ;
            rom[4811] = 8'h22 ;
            rom[4812] = 8'hf7 ;
            rom[4813] = 8'h20 ;
            rom[4814] = 8'hca ;
            rom[4815] = 8'h0d ;
            rom[4816] = 8'hf2 ;
            rom[4817] = 8'h0b ;
            rom[4818] = 8'hfb ;
            rom[4819] = 8'h23 ;
            rom[4820] = 8'h28 ;
            rom[4821] = 8'hea ;
            rom[4822] = 8'h07 ;
            rom[4823] = 8'hb2 ;
            rom[4824] = 8'hfe ;
            rom[4825] = 8'he3 ;
            rom[4826] = 8'hff ;
            rom[4827] = 8'hf4 ;
            rom[4828] = 8'h07 ;
            rom[4829] = 8'h2e ;
            rom[4830] = 8'hc8 ;
            rom[4831] = 8'hee ;
            rom[4832] = 8'h1c ;
            rom[4833] = 8'h0f ;
            rom[4834] = 8'h19 ;
            rom[4835] = 8'hbe ;
            rom[4836] = 8'h15 ;
            rom[4837] = 8'hef ;
            rom[4838] = 8'h0c ;
            rom[4839] = 8'h1d ;
            rom[4840] = 8'he5 ;
            rom[4841] = 8'hee ;
            rom[4842] = 8'hed ;
            rom[4843] = 8'hed ;
            rom[4844] = 8'hd9 ;
            rom[4845] = 8'hee ;
            rom[4846] = 8'h05 ;
            rom[4847] = 8'h28 ;
            rom[4848] = 8'hee ;
            rom[4849] = 8'hff ;
            rom[4850] = 8'h25 ;
            rom[4851] = 8'hf2 ;
            rom[4852] = 8'h08 ;
            rom[4853] = 8'hf8 ;
            rom[4854] = 8'h08 ;
            rom[4855] = 8'h02 ;
            rom[4856] = 8'he3 ;
            rom[4857] = 8'hff ;
            rom[4858] = 8'hf6 ;
            rom[4859] = 8'hea ;
            rom[4860] = 8'hdb ;
            rom[4861] = 8'hd8 ;
            rom[4862] = 8'hcf ;
            rom[4863] = 8'h0c ;
            rom[4864] = 8'hd8 ;
            rom[4865] = 8'hf2 ;
            rom[4866] = 8'hce ;
            rom[4867] = 8'h13 ;
            rom[4868] = 8'h06 ;
            rom[4869] = 8'hf6 ;
            rom[4870] = 8'he4 ;
            rom[4871] = 8'h1f ;
            rom[4872] = 8'hfe ;
            rom[4873] = 8'hcd ;
            rom[4874] = 8'hff ;
            rom[4875] = 8'hf6 ;
            rom[4876] = 8'hf6 ;
            rom[4877] = 8'he9 ;
            rom[4878] = 8'hfa ;
            rom[4879] = 8'h0d ;
            rom[4880] = 8'hf2 ;
            rom[4881] = 8'h17 ;
            rom[4882] = 8'h19 ;
            rom[4883] = 8'hf0 ;
            rom[4884] = 8'h17 ;
            rom[4885] = 8'hf2 ;
            rom[4886] = 8'h05 ;
            rom[4887] = 8'hff ;
            rom[4888] = 8'h1e ;
            rom[4889] = 8'hf9 ;
            rom[4890] = 8'h13 ;
            rom[4891] = 8'h20 ;
            rom[4892] = 8'hc9 ;
            rom[4893] = 8'h1f ;
            rom[4894] = 8'h0b ;
            rom[4895] = 8'h10 ;
            rom[4896] = 8'hff ;
            rom[4897] = 8'hc6 ;
            rom[4898] = 8'he2 ;
            rom[4899] = 8'h07 ;
            rom[4900] = 8'hfc ;
            rom[4901] = 8'he3 ;
            rom[4902] = 8'h07 ;
            rom[4903] = 8'h1c ;
            rom[4904] = 8'h1d ;
            rom[4905] = 8'hda ;
            rom[4906] = 8'hd2 ;
            rom[4907] = 8'h19 ;
            rom[4908] = 8'h06 ;
            rom[4909] = 8'h15 ;
            rom[4910] = 8'hfe ;
            rom[4911] = 8'hd9 ;
            rom[4912] = 8'h10 ;
            rom[4913] = 8'h05 ;
            rom[4914] = 8'hdc ;
            rom[4915] = 8'h02 ;
            rom[4916] = 8'he7 ;
            rom[4917] = 8'h0f ;
            rom[4918] = 8'h1e ;
            rom[4919] = 8'h15 ;
            rom[4920] = 8'hfc ;
            rom[4921] = 8'hfa ;
            rom[4922] = 8'h16 ;
            rom[4923] = 8'h11 ;
            rom[4924] = 8'hd2 ;
            rom[4925] = 8'hef ;
            rom[4926] = 8'h24 ;
            rom[4927] = 8'hf3 ;
            rom[4928] = 8'h08 ;
            rom[4929] = 8'h08 ;
            rom[4930] = 8'h0f ;
            rom[4931] = 8'hf2 ;
            rom[4932] = 8'h08 ;
            rom[4933] = 8'hfb ;
            rom[4934] = 8'hee ;
            rom[4935] = 8'h15 ;
            rom[4936] = 8'h02 ;
            rom[4937] = 8'hdf ;
            rom[4938] = 8'h01 ;
            rom[4939] = 8'h1e ;
            rom[4940] = 8'hf9 ;
            rom[4941] = 8'hc6 ;
            rom[4942] = 8'h02 ;
            rom[4943] = 8'hf3 ;
            rom[4944] = 8'hf6 ;
            rom[4945] = 8'h0d ;
            rom[4946] = 8'h0f ;
            rom[4947] = 8'he1 ;
            rom[4948] = 8'hd4 ;
            rom[4949] = 8'h0a ;
            rom[4950] = 8'hf3 ;
            rom[4951] = 8'hf5 ;
            rom[4952] = 8'h1b ;
            rom[4953] = 8'h33 ;
            rom[4954] = 8'h1a ;
            rom[4955] = 8'h04 ;
            rom[4956] = 8'h03 ;
            rom[4957] = 8'h00 ;
            rom[4958] = 8'hff ;
            rom[4959] = 8'hed ;
            rom[4960] = 8'h04 ;
            rom[4961] = 8'h24 ;
            rom[4962] = 8'h13 ;
            rom[4963] = 8'hd7 ;
            rom[4964] = 8'h05 ;
            rom[4965] = 8'he1 ;
            rom[4966] = 8'h1d ;
            rom[4967] = 8'he2 ;
            rom[4968] = 8'h16 ;
            rom[4969] = 8'h12 ;
            rom[4970] = 8'hcf ;
            rom[4971] = 8'hfa ;
            rom[4972] = 8'h03 ;
            rom[4973] = 8'h03 ;
            rom[4974] = 8'hd6 ;
            rom[4975] = 8'h04 ;
            rom[4976] = 8'h00 ;
            rom[4977] = 8'h16 ;
            rom[4978] = 8'h0b ;
            rom[4979] = 8'h04 ;
            rom[4980] = 8'h14 ;
            rom[4981] = 8'hd9 ;
            rom[4982] = 8'hf5 ;
            rom[4983] = 8'h07 ;
            rom[4984] = 8'h27 ;
            rom[4985] = 8'h15 ;
            rom[4986] = 8'h08 ;
            rom[4987] = 8'h07 ;
            rom[4988] = 8'hf9 ;
            rom[4989] = 8'hff ;
            rom[4990] = 8'hfd ;
            rom[4991] = 8'h0d ;
            rom[4992] = 8'he4 ;
            rom[4993] = 8'h0d ;
            rom[4994] = 8'h1c ;
            rom[4995] = 8'hd3 ;
            rom[4996] = 8'h06 ;
            rom[4997] = 8'h11 ;
            rom[4998] = 8'hf8 ;
            rom[4999] = 8'hdc ;
            rom[5000] = 8'h16 ;
            rom[5001] = 8'hf8 ;
            rom[5002] = 8'h02 ;
            rom[5003] = 8'hfe ;
            rom[5004] = 8'hf6 ;
            rom[5005] = 8'he4 ;
            rom[5006] = 8'h13 ;
            rom[5007] = 8'hd6 ;
            rom[5008] = 8'hce ;
            rom[5009] = 8'h1f ;
            rom[5010] = 8'h1a ;
            rom[5011] = 8'h1f ;
            rom[5012] = 8'h0b ;
            rom[5013] = 8'hfb ;
            rom[5014] = 8'h13 ;
            rom[5015] = 8'h2b ;
            rom[5016] = 8'hfc ;
            rom[5017] = 8'hee ;
            rom[5018] = 8'h12 ;
            rom[5019] = 8'h30 ;
            rom[5020] = 8'he1 ;
            rom[5021] = 8'hf7 ;
            rom[5022] = 8'h01 ;
            rom[5023] = 8'he2 ;
            rom[5024] = 8'h13 ;
            rom[5025] = 8'h0a ;
            rom[5026] = 8'h0f ;
            rom[5027] = 8'h09 ;
            rom[5028] = 8'hdf ;
            rom[5029] = 8'h0f ;
            rom[5030] = 8'hed ;
            rom[5031] = 8'hcd ;
            rom[5032] = 8'h06 ;
            rom[5033] = 8'hfc ;
            rom[5034] = 8'hef ;
            rom[5035] = 8'h04 ;
            rom[5036] = 8'h0c ;
            rom[5037] = 8'hd3 ;
            rom[5038] = 8'h00 ;
            rom[5039] = 8'he8 ;
            rom[5040] = 8'hdf ;
            rom[5041] = 8'hee ;
            rom[5042] = 8'h1a ;
            rom[5043] = 8'hdc ;
            rom[5044] = 8'h29 ;
            rom[5045] = 8'heb ;
            rom[5046] = 8'h03 ;
            rom[5047] = 8'h24 ;
            rom[5048] = 8'h03 ;
            rom[5049] = 8'h0f ;
            rom[5050] = 8'hfa ;
            rom[5051] = 8'hc9 ;
            rom[5052] = 8'h1b ;
            rom[5053] = 8'hdd ;
            rom[5054] = 8'hd8 ;
            rom[5055] = 8'he7 ;
            rom[5056] = 8'hfd ;
            rom[5057] = 8'he9 ;
            rom[5058] = 8'hd9 ;
            rom[5059] = 8'hf7 ;
            rom[5060] = 8'h11 ;
            rom[5061] = 8'h0e ;
            rom[5062] = 8'hec ;
            rom[5063] = 8'h24 ;
            rom[5064] = 8'he9 ;
            rom[5065] = 8'h0b ;
            rom[5066] = 8'h0e ;
            rom[5067] = 8'he1 ;
            rom[5068] = 8'hfb ;
            rom[5069] = 8'h15 ;
            rom[5070] = 8'hf5 ;
            rom[5071] = 8'hee ;
            rom[5072] = 8'hf9 ;
            rom[5073] = 8'h06 ;
            rom[5074] = 8'hfe ;
            rom[5075] = 8'hfb ;
            rom[5076] = 8'h19 ;
            rom[5077] = 8'hfc ;
            rom[5078] = 8'h07 ;
            rom[5079] = 8'h0b ;
            rom[5080] = 8'he2 ;
            rom[5081] = 8'h1c ;
            rom[5082] = 8'h01 ;
            rom[5083] = 8'hcd ;
            rom[5084] = 8'hfe ;
            rom[5085] = 8'hfc ;
            rom[5086] = 8'h18 ;
            rom[5087] = 8'h15 ;
            rom[5088] = 8'hf2 ;
            rom[5089] = 8'h1e ;
            rom[5090] = 8'hda ;
            rom[5091] = 8'h0f ;
            rom[5092] = 8'hd9 ;
            rom[5093] = 8'he4 ;
            rom[5094] = 8'h11 ;
            rom[5095] = 8'h02 ;
            rom[5096] = 8'h07 ;
            rom[5097] = 8'hc6 ;
            rom[5098] = 8'hce ;
            rom[5099] = 8'h13 ;
            rom[5100] = 8'hdb ;
            rom[5101] = 8'h06 ;
            rom[5102] = 8'hcd ;
            rom[5103] = 8'hf3 ;
            rom[5104] = 8'hda ;
            rom[5105] = 8'hee ;
            rom[5106] = 8'h07 ;
            rom[5107] = 8'hfb ;
            rom[5108] = 8'hf9 ;
            rom[5109] = 8'h10 ;
            rom[5110] = 8'h17 ;
            rom[5111] = 8'hf7 ;
            rom[5112] = 8'h04 ;
            rom[5113] = 8'h0e ;
            rom[5114] = 8'hf5 ;
            rom[5115] = 8'hee ;
            rom[5116] = 8'h17 ;
            rom[5117] = 8'hf4 ;
            rom[5118] = 8'h1b ;
            rom[5119] = 8'he9 ;
            rom[5120] = 8'h09 ;
            rom[5121] = 8'h06 ;
            rom[5122] = 8'hef ;
            rom[5123] = 8'h23 ;
            rom[5124] = 8'hea ;
            rom[5125] = 8'ha6 ;
            rom[5126] = 8'h0a ;
            rom[5127] = 8'he1 ;
            rom[5128] = 8'hfd ;
            rom[5129] = 8'h0b ;
            rom[5130] = 8'hef ;
            rom[5131] = 8'h11 ;
            rom[5132] = 8'h06 ;
            rom[5133] = 8'h16 ;
            rom[5134] = 8'h11 ;
            rom[5135] = 8'he6 ;
            rom[5136] = 8'h11 ;
            rom[5137] = 8'hf8 ;
            rom[5138] = 8'hf6 ;
            rom[5139] = 8'hea ;
            rom[5140] = 8'hf5 ;
            rom[5141] = 8'hff ;
            rom[5142] = 8'h04 ;
            rom[5143] = 8'h1d ;
            rom[5144] = 8'h05 ;
            rom[5145] = 8'hf9 ;
            rom[5146] = 8'he1 ;
            rom[5147] = 8'h03 ;
            rom[5148] = 8'h04 ;
            rom[5149] = 8'h1a ;
            rom[5150] = 8'hfc ;
            rom[5151] = 8'he8 ;
            rom[5152] = 8'he3 ;
            rom[5153] = 8'h02 ;
            rom[5154] = 8'hfc ;
            rom[5155] = 8'he3 ;
            rom[5156] = 8'hf2 ;
            rom[5157] = 8'he6 ;
            rom[5158] = 8'he3 ;
            rom[5159] = 8'hec ;
            rom[5160] = 8'hd4 ;
            rom[5161] = 8'he2 ;
            rom[5162] = 8'h1c ;
            rom[5163] = 8'hf8 ;
            rom[5164] = 8'hf6 ;
            rom[5165] = 8'h14 ;
            rom[5166] = 8'hd6 ;
            rom[5167] = 8'h0b ;
            rom[5168] = 8'hfd ;
            rom[5169] = 8'h10 ;
            rom[5170] = 8'hdd ;
            rom[5171] = 8'h11 ;
            rom[5172] = 8'h16 ;
            rom[5173] = 8'hf2 ;
            rom[5174] = 8'hfb ;
            rom[5175] = 8'he3 ;
            rom[5176] = 8'hf0 ;
            rom[5177] = 8'hf5 ;
            rom[5178] = 8'hf8 ;
            rom[5179] = 8'hd1 ;
            rom[5180] = 8'h0d ;
            rom[5181] = 8'hff ;
            rom[5182] = 8'hf9 ;
            rom[5183] = 8'hf3 ;
            rom[5184] = 8'h05 ;
            rom[5185] = 8'h0b ;
            rom[5186] = 8'hfd ;
            rom[5187] = 8'h01 ;
            rom[5188] = 8'h03 ;
            rom[5189] = 8'h1f ;
            rom[5190] = 8'hea ;
            rom[5191] = 8'hcc ;
            rom[5192] = 8'he7 ;
            rom[5193] = 8'h0e ;
            rom[5194] = 8'h0d ;
            rom[5195] = 8'hf6 ;
            rom[5196] = 8'he3 ;
            rom[5197] = 8'h1b ;
            rom[5198] = 8'hfd ;
            rom[5199] = 8'hec ;
            rom[5200] = 8'hf9 ;
            rom[5201] = 8'h03 ;
            rom[5202] = 8'h15 ;
            rom[5203] = 8'hf7 ;
            rom[5204] = 8'he1 ;
            rom[5205] = 8'he9 ;
            rom[5206] = 8'hdd ;
            rom[5207] = 8'hfa ;
            rom[5208] = 8'heb ;
            rom[5209] = 8'hbc ;
            rom[5210] = 8'h04 ;
            rom[5211] = 8'hd5 ;
            rom[5212] = 8'hfb ;
            rom[5213] = 8'h04 ;
            rom[5214] = 8'h22 ;
            rom[5215] = 8'hf6 ;
            rom[5216] = 8'h2e ;
            rom[5217] = 8'h14 ;
            rom[5218] = 8'hf9 ;
            rom[5219] = 8'h31 ;
            rom[5220] = 8'h00 ;
            rom[5221] = 8'h1a ;
            rom[5222] = 8'hd8 ;
            rom[5223] = 8'hf6 ;
            rom[5224] = 8'hcc ;
            rom[5225] = 8'h06 ;
            rom[5226] = 8'hf3 ;
            rom[5227] = 8'h0e ;
            rom[5228] = 8'hf2 ;
            rom[5229] = 8'h29 ;
            rom[5230] = 8'h22 ;
            rom[5231] = 8'h0a ;
            rom[5232] = 8'hfb ;
            rom[5233] = 8'hfa ;
            rom[5234] = 8'hde ;
            rom[5235] = 8'hfa ;
            rom[5236] = 8'hd6 ;
            rom[5237] = 8'h0e ;
            rom[5238] = 8'hd2 ;
            rom[5239] = 8'h02 ;
            rom[5240] = 8'hd4 ;
            rom[5241] = 8'he6 ;
            rom[5242] = 8'hdc ;
            rom[5243] = 8'hff ;
            rom[5244] = 8'hfa ;
            rom[5245] = 8'he5 ;
            rom[5246] = 8'h05 ;
            rom[5247] = 8'h07 ;
            rom[5248] = 8'hda ;
            rom[5249] = 8'h0a ;
            rom[5250] = 8'h0e ;
            rom[5251] = 8'hfa ;
            rom[5252] = 8'h08 ;
            rom[5253] = 8'hee ;
            rom[5254] = 8'hf9 ;
            rom[5255] = 8'hfd ;
            rom[5256] = 8'hd2 ;
            rom[5257] = 8'h21 ;
            rom[5258] = 8'h0a ;
            rom[5259] = 8'hef ;
            rom[5260] = 8'hd9 ;
            rom[5261] = 8'h2f ;
            rom[5262] = 8'hfb ;
            rom[5263] = 8'h05 ;
            rom[5264] = 8'he6 ;
            rom[5265] = 8'h22 ;
            rom[5266] = 8'he2 ;
            rom[5267] = 8'hd4 ;
            rom[5268] = 8'h0a ;
            rom[5269] = 8'h24 ;
            rom[5270] = 8'hef ;
            rom[5271] = 8'h07 ;
            rom[5272] = 8'h20 ;
            rom[5273] = 8'h28 ;
            rom[5274] = 8'h0c ;
            rom[5275] = 8'h20 ;
            rom[5276] = 8'h13 ;
            rom[5277] = 8'h16 ;
            rom[5278] = 8'h02 ;
            rom[5279] = 8'hf1 ;
            rom[5280] = 8'hff ;
            rom[5281] = 8'h14 ;
            rom[5282] = 8'h0c ;
            rom[5283] = 8'h11 ;
            rom[5284] = 8'hf2 ;
            rom[5285] = 8'hf2 ;
            rom[5286] = 8'hf7 ;
            rom[5287] = 8'he7 ;
            rom[5288] = 8'hec ;
            rom[5289] = 8'hfb ;
            rom[5290] = 8'hfb ;
            rom[5291] = 8'hf0 ;
            rom[5292] = 8'hfd ;
            rom[5293] = 8'hb8 ;
            rom[5294] = 8'h03 ;
            rom[5295] = 8'hd4 ;
            rom[5296] = 8'he9 ;
            rom[5297] = 8'he3 ;
            rom[5298] = 8'hf3 ;
            rom[5299] = 8'hdb ;
            rom[5300] = 8'h14 ;
            rom[5301] = 8'h0e ;
            rom[5302] = 8'hf9 ;
            rom[5303] = 8'hfc ;
            rom[5304] = 8'h28 ;
            rom[5305] = 8'hda ;
            rom[5306] = 8'hf6 ;
            rom[5307] = 8'hef ;
            rom[5308] = 8'h06 ;
            rom[5309] = 8'hd3 ;
            rom[5310] = 8'h0b ;
            rom[5311] = 8'hf3 ;
            rom[5312] = 8'hf3 ;
            rom[5313] = 8'h17 ;
            rom[5314] = 8'hf7 ;
            rom[5315] = 8'h13 ;
            rom[5316] = 8'hf5 ;
            rom[5317] = 8'hde ;
            rom[5318] = 8'h02 ;
            rom[5319] = 8'h0e ;
            rom[5320] = 8'hec ;
            rom[5321] = 8'h03 ;
            rom[5322] = 8'h0c ;
            rom[5323] = 8'h0f ;
            rom[5324] = 8'h02 ;
            rom[5325] = 8'hfb ;
            rom[5326] = 8'h19 ;
            rom[5327] = 8'h07 ;
            rom[5328] = 8'hda ;
            rom[5329] = 8'h0b ;
            rom[5330] = 8'hf0 ;
            rom[5331] = 8'h1a ;
            rom[5332] = 8'h13 ;
            rom[5333] = 8'h09 ;
            rom[5334] = 8'h14 ;
            rom[5335] = 8'hef ;
            rom[5336] = 8'h08 ;
            rom[5337] = 8'h14 ;
            rom[5338] = 8'hd7 ;
            rom[5339] = 8'hf3 ;
            rom[5340] = 8'h08 ;
            rom[5341] = 8'h2e ;
            rom[5342] = 8'h06 ;
            rom[5343] = 8'he3 ;
            rom[5344] = 8'hea ;
            rom[5345] = 8'hfd ;
            rom[5346] = 8'h11 ;
            rom[5347] = 8'hb4 ;
            rom[5348] = 8'h01 ;
            rom[5349] = 8'h9d ;
            rom[5350] = 8'he0 ;
            rom[5351] = 8'h23 ;
            rom[5352] = 8'h0b ;
            rom[5353] = 8'h28 ;
            rom[5354] = 8'hc0 ;
            rom[5355] = 8'hf7 ;
            rom[5356] = 8'hf3 ;
            rom[5357] = 8'hde ;
            rom[5358] = 8'hed ;
            rom[5359] = 8'h11 ;
            rom[5360] = 8'hf1 ;
            rom[5361] = 8'h09 ;
            rom[5362] = 8'h06 ;
            rom[5363] = 8'h2b ;
            rom[5364] = 8'he7 ;
            rom[5365] = 8'hda ;
            rom[5366] = 8'h12 ;
            rom[5367] = 8'h04 ;
            rom[5368] = 8'hea ;
            rom[5369] = 8'h3e ;
            rom[5370] = 8'hf4 ;
            rom[5371] = 8'he1 ;
            rom[5372] = 8'hfb ;
            rom[5373] = 8'h15 ;
            rom[5374] = 8'hf4 ;
            rom[5375] = 8'h24 ;
            rom[5376] = 8'hd1 ;
            rom[5377] = 8'hf1 ;
            rom[5378] = 8'heb ;
            rom[5379] = 8'hfd ;
            rom[5380] = 8'h0a ;
            rom[5381] = 8'h1a ;
            rom[5382] = 8'hed ;
            rom[5383] = 8'h22 ;
            rom[5384] = 8'hf8 ;
            rom[5385] = 8'he5 ;
            rom[5386] = 8'h0d ;
            rom[5387] = 8'hd3 ;
            rom[5388] = 8'h15 ;
            rom[5389] = 8'hff ;
            rom[5390] = 8'h14 ;
            rom[5391] = 8'h13 ;
            rom[5392] = 8'h07 ;
            rom[5393] = 8'hfe ;
            rom[5394] = 8'h03 ;
            rom[5395] = 8'h07 ;
            rom[5396] = 8'heb ;
            rom[5397] = 8'he8 ;
            rom[5398] = 8'hfe ;
            rom[5399] = 8'h2e ;
            rom[5400] = 8'h08 ;
            rom[5401] = 8'hf7 ;
            rom[5402] = 8'h0e ;
            rom[5403] = 8'hf3 ;
            rom[5404] = 8'h04 ;
            rom[5405] = 8'h12 ;
            rom[5406] = 8'hdf ;
            rom[5407] = 8'hcd ;
            rom[5408] = 8'h03 ;
            rom[5409] = 8'hfa ;
            rom[5410] = 8'hf6 ;
            rom[5411] = 8'hf3 ;
            rom[5412] = 8'hee ;
            rom[5413] = 8'h01 ;
            rom[5414] = 8'h05 ;
            rom[5415] = 8'h29 ;
            rom[5416] = 8'hfb ;
            rom[5417] = 8'he1 ;
            rom[5418] = 8'h0f ;
            rom[5419] = 8'h09 ;
            rom[5420] = 8'hf3 ;
            rom[5421] = 8'h0c ;
            rom[5422] = 8'h15 ;
            rom[5423] = 8'he4 ;
            rom[5424] = 8'he2 ;
            rom[5425] = 8'h0e ;
            rom[5426] = 8'h08 ;
            rom[5427] = 8'hec ;
            rom[5428] = 8'hca ;
            rom[5429] = 8'h05 ;
            rom[5430] = 8'h2c ;
            rom[5431] = 8'h05 ;
            rom[5432] = 8'h01 ;
            rom[5433] = 8'hfe ;
            rom[5434] = 8'h08 ;
            rom[5435] = 8'hd5 ;
            rom[5436] = 8'he2 ;
            rom[5437] = 8'hf9 ;
            rom[5438] = 8'hf9 ;
            rom[5439] = 8'h24 ;
            rom[5440] = 8'h15 ;
            rom[5441] = 8'he8 ;
            rom[5442] = 8'h0d ;
            rom[5443] = 8'hfa ;
            rom[5444] = 8'hec ;
            rom[5445] = 8'hee ;
            rom[5446] = 8'h10 ;
            rom[5447] = 8'hf4 ;
            rom[5448] = 8'h1c ;
            rom[5449] = 8'ha2 ;
            rom[5450] = 8'hfd ;
            rom[5451] = 8'hf7 ;
            rom[5452] = 8'hff ;
            rom[5453] = 8'h0d ;
            rom[5454] = 8'hc4 ;
            rom[5455] = 8'h04 ;
            rom[5456] = 8'h30 ;
            rom[5457] = 8'hfa ;
            rom[5458] = 8'h03 ;
            rom[5459] = 8'h1a ;
            rom[5460] = 8'hfe ;
            rom[5461] = 8'hdd ;
            rom[5462] = 8'h16 ;
            rom[5463] = 8'hdc ;
            rom[5464] = 8'h02 ;
            rom[5465] = 8'hf0 ;
            rom[5466] = 8'h14 ;
            rom[5467] = 8'hff ;
            rom[5468] = 8'he9 ;
            rom[5469] = 8'h08 ;
            rom[5470] = 8'he6 ;
            rom[5471] = 8'h01 ;
            rom[5472] = 8'h01 ;
            rom[5473] = 8'hf8 ;
            rom[5474] = 8'hfd ;
            rom[5475] = 8'hdb ;
            rom[5476] = 8'h07 ;
            rom[5477] = 8'hd9 ;
            rom[5478] = 8'h2e ;
            rom[5479] = 8'h06 ;
            rom[5480] = 8'hd1 ;
            rom[5481] = 8'hd0 ;
            rom[5482] = 8'hfc ;
            rom[5483] = 8'h0b ;
            rom[5484] = 8'he7 ;
            rom[5485] = 8'h05 ;
            rom[5486] = 8'he3 ;
            rom[5487] = 8'hf4 ;
            rom[5488] = 8'h22 ;
            rom[5489] = 8'hed ;
            rom[5490] = 8'h39 ;
            rom[5491] = 8'hf2 ;
            rom[5492] = 8'hd2 ;
            rom[5493] = 8'hea ;
            rom[5494] = 8'he9 ;
            rom[5495] = 8'hf8 ;
            rom[5496] = 8'hd3 ;
            rom[5497] = 8'h0c ;
            rom[5498] = 8'h22 ;
            rom[5499] = 8'h07 ;
            rom[5500] = 8'hf4 ;
            rom[5501] = 8'he1 ;
            rom[5502] = 8'h13 ;
            rom[5503] = 8'h0a ;
            rom[5504] = 8'h09 ;
            rom[5505] = 8'h23 ;
            rom[5506] = 8'he8 ;
            rom[5507] = 8'h0e ;
            rom[5508] = 8'he6 ;
            rom[5509] = 8'hcd ;
            rom[5510] = 8'hfd ;
            rom[5511] = 8'hde ;
            rom[5512] = 8'hfd ;
            rom[5513] = 8'h0d ;
            rom[5514] = 8'hda ;
            rom[5515] = 8'hff ;
            rom[5516] = 8'hff ;
            rom[5517] = 8'h08 ;
            rom[5518] = 8'hf9 ;
            rom[5519] = 8'h16 ;
            rom[5520] = 8'h0c ;
            rom[5521] = 8'he9 ;
            rom[5522] = 8'hb3 ;
            rom[5523] = 8'he0 ;
            rom[5524] = 8'h22 ;
            rom[5525] = 8'h2b ;
            rom[5526] = 8'h10 ;
            rom[5527] = 8'hf6 ;
            rom[5528] = 8'hf4 ;
            rom[5529] = 8'hfe ;
            rom[5530] = 8'hdf ;
            rom[5531] = 8'hfc ;
            rom[5532] = 8'hf4 ;
            rom[5533] = 8'hfe ;
            rom[5534] = 8'h1b ;
            rom[5535] = 8'hd9 ;
            rom[5536] = 8'h09 ;
            rom[5537] = 8'hf7 ;
            rom[5538] = 8'h0e ;
            rom[5539] = 8'he7 ;
            rom[5540] = 8'h09 ;
            rom[5541] = 8'h13 ;
            rom[5542] = 8'hf0 ;
            rom[5543] = 8'h15 ;
            rom[5544] = 8'hea ;
            rom[5545] = 8'hfd ;
            rom[5546] = 8'h0a ;
            rom[5547] = 8'hec ;
            rom[5548] = 8'h0d ;
            rom[5549] = 8'hef ;
            rom[5550] = 8'hfa ;
            rom[5551] = 8'hf5 ;
            rom[5552] = 8'he4 ;
            rom[5553] = 8'h02 ;
            rom[5554] = 8'hd0 ;
            rom[5555] = 8'hf2 ;
            rom[5556] = 8'h0e ;
            rom[5557] = 8'hf7 ;
            rom[5558] = 8'hc5 ;
            rom[5559] = 8'hd5 ;
            rom[5560] = 8'hfa ;
            rom[5561] = 8'h01 ;
            rom[5562] = 8'hc7 ;
            rom[5563] = 8'h01 ;
            rom[5564] = 8'hf6 ;
            rom[5565] = 8'hf9 ;
            rom[5566] = 8'ha9 ;
            rom[5567] = 8'he5 ;
            rom[5568] = 8'hfc ;
            rom[5569] = 8'h09 ;
            rom[5570] = 8'h20 ;
            rom[5571] = 8'he6 ;
            rom[5572] = 8'hed ;
            rom[5573] = 8'he6 ;
            rom[5574] = 8'h04 ;
            rom[5575] = 8'hd7 ;
            rom[5576] = 8'hfd ;
            rom[5577] = 8'he8 ;
            rom[5578] = 8'h12 ;
            rom[5579] = 8'h06 ;
            rom[5580] = 8'hef ;
            rom[5581] = 8'h15 ;
            rom[5582] = 8'hf2 ;
            rom[5583] = 8'h02 ;
            rom[5584] = 8'h12 ;
            rom[5585] = 8'h19 ;
            rom[5586] = 8'he2 ;
            rom[5587] = 8'h0b ;
            rom[5588] = 8'he0 ;
            rom[5589] = 8'hf5 ;
            rom[5590] = 8'hed ;
            rom[5591] = 8'hf5 ;
            rom[5592] = 8'hf5 ;
            rom[5593] = 8'h06 ;
            rom[5594] = 8'hfb ;
            rom[5595] = 8'hfc ;
            rom[5596] = 8'hfa ;
            rom[5597] = 8'h0e ;
            rom[5598] = 8'hf3 ;
            rom[5599] = 8'hf3 ;
            rom[5600] = 8'he5 ;
            rom[5601] = 8'hfb ;
            rom[5602] = 8'hcb ;
            rom[5603] = 8'hfd ;
            rom[5604] = 8'h0b ;
            rom[5605] = 8'hff ;
            rom[5606] = 8'hdc ;
            rom[5607] = 8'h04 ;
            rom[5608] = 8'hde ;
            rom[5609] = 8'hf6 ;
            rom[5610] = 8'h08 ;
            rom[5611] = 8'hdb ;
            rom[5612] = 8'he5 ;
            rom[5613] = 8'hd9 ;
            rom[5614] = 8'hee ;
            rom[5615] = 8'h2c ;
            rom[5616] = 8'hfd ;
            rom[5617] = 8'hfb ;
            rom[5618] = 8'h15 ;
            rom[5619] = 8'he4 ;
            rom[5620] = 8'hf8 ;
            rom[5621] = 8'hf3 ;
            rom[5622] = 8'hf6 ;
            rom[5623] = 8'he5 ;
            rom[5624] = 8'hd7 ;
            rom[5625] = 8'h08 ;
            rom[5626] = 8'hfd ;
            rom[5627] = 8'hd4 ;
            rom[5628] = 8'h04 ;
            rom[5629] = 8'hab ;
            rom[5630] = 8'hf0 ;
            rom[5631] = 8'h02 ;
            rom[5632] = 8'hda ;
            rom[5633] = 8'hdf ;
            rom[5634] = 8'h05 ;
            rom[5635] = 8'hfa ;
            rom[5636] = 8'he9 ;
            rom[5637] = 8'hfd ;
            rom[5638] = 8'hf6 ;
            rom[5639] = 8'hee ;
            rom[5640] = 8'h00 ;
            rom[5641] = 8'hb9 ;
            rom[5642] = 8'hf9 ;
            rom[5643] = 8'hf4 ;
            rom[5644] = 8'h0c ;
            rom[5645] = 8'hee ;
            rom[5646] = 8'h04 ;
            rom[5647] = 8'h0b ;
            rom[5648] = 8'h00 ;
            rom[5649] = 8'h06 ;
            rom[5650] = 8'he6 ;
            rom[5651] = 8'hf6 ;
            rom[5652] = 8'he6 ;
            rom[5653] = 8'heb ;
            rom[5654] = 8'hf7 ;
            rom[5655] = 8'hdc ;
            rom[5656] = 8'hd5 ;
            rom[5657] = 8'h09 ;
            rom[5658] = 8'hfa ;
            rom[5659] = 8'hb3 ;
            rom[5660] = 8'h1c ;
            rom[5661] = 8'hdb ;
            rom[5662] = 8'h0d ;
            rom[5663] = 8'hf3 ;
            rom[5664] = 8'h06 ;
            rom[5665] = 8'h17 ;
            rom[5666] = 8'hf8 ;
            rom[5667] = 8'hec ;
            rom[5668] = 8'h1d ;
            rom[5669] = 8'hfe ;
            rom[5670] = 8'hf6 ;
            rom[5671] = 8'he4 ;
            rom[5672] = 8'h0b ;
            rom[5673] = 8'heb ;
            rom[5674] = 8'h1f ;
            rom[5675] = 8'hf1 ;
            rom[5676] = 8'hcf ;
            rom[5677] = 8'hf2 ;
            rom[5678] = 8'he2 ;
            rom[5679] = 8'h02 ;
            rom[5680] = 8'hf4 ;
            rom[5681] = 8'hda ;
            rom[5682] = 8'he5 ;
            rom[5683] = 8'h09 ;
            rom[5684] = 8'hf8 ;
            rom[5685] = 8'hf0 ;
            rom[5686] = 8'hfd ;
            rom[5687] = 8'h19 ;
            rom[5688] = 8'hc6 ;
            rom[5689] = 8'h1f ;
            rom[5690] = 8'hb7 ;
            rom[5691] = 8'hf4 ;
            rom[5692] = 8'hea ;
            rom[5693] = 8'h1a ;
            rom[5694] = 8'hf1 ;
            rom[5695] = 8'h06 ;
            rom[5696] = 8'h12 ;
            rom[5697] = 8'hf1 ;
            rom[5698] = 8'h33 ;
            rom[5699] = 8'h01 ;
            rom[5700] = 8'h10 ;
            rom[5701] = 8'hfa ;
            rom[5702] = 8'hff ;
            rom[5703] = 8'hf0 ;
            rom[5704] = 8'h09 ;
            rom[5705] = 8'hce ;
            rom[5706] = 8'hfb ;
            rom[5707] = 8'h08 ;
            rom[5708] = 8'hca ;
            rom[5709] = 8'h01 ;
            rom[5710] = 8'he9 ;
            rom[5711] = 8'h04 ;
            rom[5712] = 8'hec ;
            rom[5713] = 8'hea ;
            rom[5714] = 8'h03 ;
            rom[5715] = 8'hf0 ;
            rom[5716] = 8'h0c ;
            rom[5717] = 8'hf6 ;
            rom[5718] = 8'hf2 ;
            rom[5719] = 8'h1f ;
            rom[5720] = 8'hf4 ;
            rom[5721] = 8'h2b ;
            rom[5722] = 8'hf0 ;
            rom[5723] = 8'h18 ;
            rom[5724] = 8'hfc ;
            rom[5725] = 8'hf5 ;
            rom[5726] = 8'h06 ;
            rom[5727] = 8'h07 ;
            rom[5728] = 8'hcb ;
            rom[5729] = 8'hed ;
            rom[5730] = 8'hc6 ;
            rom[5731] = 8'hfd ;
            rom[5732] = 8'hed ;
            rom[5733] = 8'he1 ;
            rom[5734] = 8'h04 ;
            rom[5735] = 8'hfe ;
            rom[5736] = 8'hfa ;
            rom[5737] = 8'hfc ;
            rom[5738] = 8'hfe ;
            rom[5739] = 8'he4 ;
            rom[5740] = 8'h09 ;
            rom[5741] = 8'h2a ;
            rom[5742] = 8'h02 ;
            rom[5743] = 8'h11 ;
            rom[5744] = 8'h11 ;
            rom[5745] = 8'hf0 ;
            rom[5746] = 8'h2c ;
            rom[5747] = 8'hf1 ;
            rom[5748] = 8'he4 ;
            rom[5749] = 8'h04 ;
            rom[5750] = 8'h10 ;
            rom[5751] = 8'h0f ;
            rom[5752] = 8'h06 ;
            rom[5753] = 8'h13 ;
            rom[5754] = 8'hdb ;
            rom[5755] = 8'hf4 ;
            rom[5756] = 8'hff ;
            rom[5757] = 8'hfd ;
            rom[5758] = 8'hd0 ;
            rom[5759] = 8'hfd ;
            rom[5760] = 8'h0e ;
            rom[5761] = 8'hf1 ;
            rom[5762] = 8'he4 ;
            rom[5763] = 8'h18 ;
            rom[5764] = 8'hfc ;
            rom[5765] = 8'hde ;
            rom[5766] = 8'h1c ;
            rom[5767] = 8'hf7 ;
            rom[5768] = 8'h1c ;
            rom[5769] = 8'hec ;
            rom[5770] = 8'he1 ;
            rom[5771] = 8'h04 ;
            rom[5772] = 8'hd7 ;
            rom[5773] = 8'h18 ;
            rom[5774] = 8'hf1 ;
            rom[5775] = 8'h11 ;
            rom[5776] = 8'hfd ;
            rom[5777] = 8'hec ;
            rom[5778] = 8'hf3 ;
            rom[5779] = 8'h03 ;
            rom[5780] = 8'hfd ;
            rom[5781] = 8'hd2 ;
            rom[5782] = 8'hdf ;
            rom[5783] = 8'h0e ;
            rom[5784] = 8'he9 ;
            rom[5785] = 8'hf4 ;
            rom[5786] = 8'hf4 ;
            rom[5787] = 8'he3 ;
            rom[5788] = 8'h03 ;
            rom[5789] = 8'h00 ;
            rom[5790] = 8'heb ;
            rom[5791] = 8'hf4 ;
            rom[5792] = 8'h20 ;
            rom[5793] = 8'h1d ;
            rom[5794] = 8'he6 ;
            rom[5795] = 8'hee ;
            rom[5796] = 8'hee ;
            rom[5797] = 8'h10 ;
            rom[5798] = 8'he9 ;
            rom[5799] = 8'h0a ;
            rom[5800] = 8'hf1 ;
            rom[5801] = 8'hf0 ;
            rom[5802] = 8'h32 ;
            rom[5803] = 8'hdf ;
            rom[5804] = 8'he5 ;
            rom[5805] = 8'h05 ;
            rom[5806] = 8'hdb ;
            rom[5807] = 8'hfc ;
            rom[5808] = 8'hfd ;
            rom[5809] = 8'hf4 ;
            rom[5810] = 8'he3 ;
            rom[5811] = 8'hf6 ;
            rom[5812] = 8'h04 ;
            rom[5813] = 8'hfa ;
            rom[5814] = 8'he5 ;
            rom[5815] = 8'h1a ;
            rom[5816] = 8'he6 ;
            rom[5817] = 8'h24 ;
            rom[5818] = 8'hdf ;
            rom[5819] = 8'he1 ;
            rom[5820] = 8'h07 ;
            rom[5821] = 8'h07 ;
            rom[5822] = 8'he4 ;
            rom[5823] = 8'he5 ;
            rom[5824] = 8'hf8 ;
            rom[5825] = 8'hfa ;
            rom[5826] = 8'he0 ;
            rom[5827] = 8'h01 ;
            rom[5828] = 8'hf1 ;
            rom[5829] = 8'h11 ;
            rom[5830] = 8'hf9 ;
            rom[5831] = 8'hd4 ;
            rom[5832] = 8'hf1 ;
            rom[5833] = 8'h1b ;
            rom[5834] = 8'hf4 ;
            rom[5835] = 8'h04 ;
            rom[5836] = 8'hfe ;
            rom[5837] = 8'h2f ;
            rom[5838] = 8'h12 ;
            rom[5839] = 8'h13 ;
            rom[5840] = 8'hf3 ;
            rom[5841] = 8'h00 ;
            rom[5842] = 8'he1 ;
            rom[5843] = 8'h02 ;
            rom[5844] = 8'hf2 ;
            rom[5845] = 8'hb8 ;
            rom[5846] = 8'h18 ;
            rom[5847] = 8'hf5 ;
            rom[5848] = 8'hfb ;
            rom[5849] = 8'h0f ;
            rom[5850] = 8'h1b ;
            rom[5851] = 8'hfb ;
            rom[5852] = 8'h02 ;
            rom[5853] = 8'hd6 ;
            rom[5854] = 8'hef ;
            rom[5855] = 8'hfc ;
            rom[5856] = 8'h0c ;
            rom[5857] = 8'hfc ;
            rom[5858] = 8'hd5 ;
            rom[5859] = 8'hf0 ;
            rom[5860] = 8'hed ;
            rom[5861] = 8'hfd ;
            rom[5862] = 8'hf8 ;
            rom[5863] = 8'hf3 ;
            rom[5864] = 8'hf0 ;
            rom[5865] = 8'hce ;
            rom[5866] = 8'hd0 ;
            rom[5867] = 8'h12 ;
            rom[5868] = 8'hf0 ;
            rom[5869] = 8'hdb ;
            rom[5870] = 8'he9 ;
            rom[5871] = 8'h1b ;
            rom[5872] = 8'h0c ;
            rom[5873] = 8'hed ;
            rom[5874] = 8'hff ;
            rom[5875] = 8'hde ;
            rom[5876] = 8'he9 ;
            rom[5877] = 8'h08 ;
            rom[5878] = 8'hea ;
            rom[5879] = 8'hcd ;
            rom[5880] = 8'hf6 ;
            rom[5881] = 8'he8 ;
            rom[5882] = 8'hdb ;
            rom[5883] = 8'h08 ;
            rom[5884] = 8'h0f ;
            rom[5885] = 8'hbd ;
            rom[5886] = 8'hfc ;
            rom[5887] = 8'hf6 ;
            rom[5888] = 8'h18 ;
            rom[5889] = 8'h00 ;
            rom[5890] = 8'hec ;
            rom[5891] = 8'he1 ;
            rom[5892] = 8'he8 ;
            rom[5893] = 8'hca ;
            rom[5894] = 8'h0f ;
            rom[5895] = 8'he3 ;
            rom[5896] = 8'hf2 ;
            rom[5897] = 8'h0f ;
            rom[5898] = 8'h00 ;
            rom[5899] = 8'h1a ;
            rom[5900] = 8'hee ;
            rom[5901] = 8'he5 ;
            rom[5902] = 8'he2 ;
            rom[5903] = 8'he3 ;
            rom[5904] = 8'hd4 ;
            rom[5905] = 8'h25 ;
            rom[5906] = 8'h04 ;
            rom[5907] = 8'hf1 ;
            rom[5908] = 8'h18 ;
            rom[5909] = 8'hea ;
            rom[5910] = 8'hd2 ;
            rom[5911] = 8'he5 ;
            rom[5912] = 8'hc6 ;
            rom[5913] = 8'h1a ;
            rom[5914] = 8'hf2 ;
            rom[5915] = 8'hd1 ;
            rom[5916] = 8'hf0 ;
            rom[5917] = 8'h15 ;
            rom[5918] = 8'h1c ;
            rom[5919] = 8'h18 ;
            rom[5920] = 8'hf4 ;
            rom[5921] = 8'hea ;
            rom[5922] = 8'h1b ;
            rom[5923] = 8'h1a ;
            rom[5924] = 8'hfd ;
            rom[5925] = 8'hef ;
            rom[5926] = 8'hf8 ;
            rom[5927] = 8'h12 ;
            rom[5928] = 8'h05 ;
            rom[5929] = 8'h03 ;
            rom[5930] = 8'hfc ;
            rom[5931] = 8'hec ;
            rom[5932] = 8'h10 ;
            rom[5933] = 8'h0a ;
            rom[5934] = 8'h15 ;
            rom[5935] = 8'hf6 ;
            rom[5936] = 8'h16 ;
            rom[5937] = 8'hfb ;
            rom[5938] = 8'hd4 ;
            rom[5939] = 8'h04 ;
            rom[5940] = 8'h07 ;
            rom[5941] = 8'he6 ;
            rom[5942] = 8'h02 ;
            rom[5943] = 8'h03 ;
            rom[5944] = 8'h0a ;
            rom[5945] = 8'h08 ;
            rom[5946] = 8'h17 ;
            rom[5947] = 8'hf8 ;
            rom[5948] = 8'h03 ;
            rom[5949] = 8'he8 ;
            rom[5950] = 8'h0d ;
            rom[5951] = 8'h07 ;
            rom[5952] = 8'hce ;
            rom[5953] = 8'hf9 ;
            rom[5954] = 8'h0d ;
            rom[5955] = 8'hdd ;
            rom[5956] = 8'hf0 ;
            rom[5957] = 8'h20 ;
            rom[5958] = 8'he3 ;
            rom[5959] = 8'h00 ;
            rom[5960] = 8'h0c ;
            rom[5961] = 8'h1c ;
            rom[5962] = 8'hf1 ;
            rom[5963] = 8'he6 ;
            rom[5964] = 8'hf9 ;
            rom[5965] = 8'hea ;
            rom[5966] = 8'h16 ;
            rom[5967] = 8'he9 ;
            rom[5968] = 8'h05 ;
            rom[5969] = 8'hf0 ;
            rom[5970] = 8'hde ;
            rom[5971] = 8'hfd ;
            rom[5972] = 8'hfe ;
            rom[5973] = 8'hf7 ;
            rom[5974] = 8'hdc ;
            rom[5975] = 8'h0f ;
            rom[5976] = 8'hef ;
            rom[5977] = 8'heb ;
            rom[5978] = 8'h14 ;
            rom[5979] = 8'he2 ;
            rom[5980] = 8'hbf ;
            rom[5981] = 8'hf0 ;
            rom[5982] = 8'h06 ;
            rom[5983] = 8'h0d ;
            rom[5984] = 8'hf6 ;
            rom[5985] = 8'hdc ;
            rom[5986] = 8'hee ;
            rom[5987] = 8'hf3 ;
            rom[5988] = 8'h15 ;
            rom[5989] = 8'h10 ;
            rom[5990] = 8'h0e ;
            rom[5991] = 8'hf8 ;
            rom[5992] = 8'hea ;
            rom[5993] = 8'h01 ;
            rom[5994] = 8'h0b ;
            rom[5995] = 8'he6 ;
            rom[5996] = 8'h00 ;
            rom[5997] = 8'h09 ;
            rom[5998] = 8'h2b ;
            rom[5999] = 8'hc7 ;
            rom[6000] = 8'hc2 ;
            rom[6001] = 8'hc7 ;
            rom[6002] = 8'hfb ;
            rom[6003] = 8'hdf ;
            rom[6004] = 8'h22 ;
            rom[6005] = 8'h1d ;
            rom[6006] = 8'hc9 ;
            rom[6007] = 8'he5 ;
            rom[6008] = 8'he3 ;
            rom[6009] = 8'hc8 ;
            rom[6010] = 8'hd5 ;
            rom[6011] = 8'h0e ;
            rom[6012] = 8'h04 ;
            rom[6013] = 8'hee ;
            rom[6014] = 8'h10 ;
            rom[6015] = 8'hbb ;
            rom[6016] = 8'hee ;
            rom[6017] = 8'he7 ;
            rom[6018] = 8'hcf ;
            rom[6019] = 8'hdc ;
            rom[6020] = 8'hdf ;
            rom[6021] = 8'hec ;
            rom[6022] = 8'hf7 ;
            rom[6023] = 8'h3a ;
            rom[6024] = 8'hdd ;
            rom[6025] = 8'h0a ;
            rom[6026] = 8'hee ;
            rom[6027] = 8'hdc ;
            rom[6028] = 8'he1 ;
            rom[6029] = 8'hf6 ;
            rom[6030] = 8'hfb ;
            rom[6031] = 8'hc0 ;
            rom[6032] = 8'h07 ;
            rom[6033] = 8'hd5 ;
            rom[6034] = 8'h14 ;
            rom[6035] = 8'h08 ;
            rom[6036] = 8'hf0 ;
            rom[6037] = 8'hf3 ;
            rom[6038] = 8'h09 ;
            rom[6039] = 8'h18 ;
            rom[6040] = 8'hf3 ;
            rom[6041] = 8'hf8 ;
            rom[6042] = 8'h13 ;
            rom[6043] = 8'hf0 ;
            rom[6044] = 8'h03 ;
            rom[6045] = 8'hf7 ;
            rom[6046] = 8'h25 ;
            rom[6047] = 8'h19 ;
            rom[6048] = 8'h2a ;
            rom[6049] = 8'h3b ;
            rom[6050] = 8'h19 ;
            rom[6051] = 8'h02 ;
            rom[6052] = 8'hf6 ;
            rom[6053] = 8'hf7 ;
            rom[6054] = 8'h19 ;
            rom[6055] = 8'hd4 ;
            rom[6056] = 8'hee ;
            rom[6057] = 8'hcf ;
            rom[6058] = 8'hed ;
            rom[6059] = 8'h05 ;
            rom[6060] = 8'h01 ;
            rom[6061] = 8'hec ;
            rom[6062] = 8'hc7 ;
            rom[6063] = 8'hf6 ;
            rom[6064] = 8'h12 ;
            rom[6065] = 8'hd2 ;
            rom[6066] = 8'h12 ;
            rom[6067] = 8'hfa ;
            rom[6068] = 8'hd4 ;
            rom[6069] = 8'h00 ;
            rom[6070] = 8'h18 ;
            rom[6071] = 8'h11 ;
            rom[6072] = 8'hf4 ;
            rom[6073] = 8'hf9 ;
            rom[6074] = 8'h1f ;
            rom[6075] = 8'hf9 ;
            rom[6076] = 8'hc6 ;
            rom[6077] = 8'h09 ;
            rom[6078] = 8'h05 ;
            rom[6079] = 8'h05 ;
            rom[6080] = 8'h20 ;
            rom[6081] = 8'hf5 ;
            rom[6082] = 8'h04 ;
            rom[6083] = 8'hc4 ;
            rom[6084] = 8'hfc ;
            rom[6085] = 8'h09 ;
            rom[6086] = 8'hf8 ;
            rom[6087] = 8'hd1 ;
            rom[6088] = 8'hfd ;
            rom[6089] = 8'he6 ;
            rom[6090] = 8'hfd ;
            rom[6091] = 8'h0c ;
            rom[6092] = 8'h0c ;
            rom[6093] = 8'hfe ;
            rom[6094] = 8'hde ;
            rom[6095] = 8'h20 ;
            rom[6096] = 8'h22 ;
            rom[6097] = 8'he2 ;
            rom[6098] = 8'h1e ;
            rom[6099] = 8'he3 ;
            rom[6100] = 8'h08 ;
            rom[6101] = 8'hef ;
            rom[6102] = 8'he4 ;
            rom[6103] = 8'hfa ;
            rom[6104] = 8'hf4 ;
            rom[6105] = 8'h15 ;
            rom[6106] = 8'h0d ;
            rom[6107] = 8'hf9 ;
            rom[6108] = 8'h21 ;
            rom[6109] = 8'hf8 ;
            rom[6110] = 8'hf8 ;
            rom[6111] = 8'h0b ;
            rom[6112] = 8'h04 ;
            rom[6113] = 8'hfd ;
            rom[6114] = 8'h00 ;
            rom[6115] = 8'h09 ;
            rom[6116] = 8'he2 ;
            rom[6117] = 8'h0c ;
            rom[6118] = 8'h2c ;
            rom[6119] = 8'hef ;
            rom[6120] = 8'h09 ;
            rom[6121] = 8'hec ;
            rom[6122] = 8'h1d ;
            rom[6123] = 8'h16 ;
            rom[6124] = 8'h0a ;
            rom[6125] = 8'h36 ;
            rom[6126] = 8'hf0 ;
            rom[6127] = 8'h15 ;
            rom[6128] = 8'h1e ;
            rom[6129] = 8'hf1 ;
            rom[6130] = 8'hf7 ;
            rom[6131] = 8'hd9 ;
            rom[6132] = 8'h0b ;
            rom[6133] = 8'hfb ;
            rom[6134] = 8'h01 ;
            rom[6135] = 8'h1f ;
            rom[6136] = 8'hf4 ;
            rom[6137] = 8'h0b ;
            rom[6138] = 8'hf9 ;
            rom[6139] = 8'h13 ;
            rom[6140] = 8'hcc ;
            rom[6141] = 8'h38 ;
            rom[6142] = 8'h0e ;
            rom[6143] = 8'h0d ;
            rom[6144] = 8'he0 ;
            rom[6145] = 8'hff ;
            rom[6146] = 8'hfb ;
            rom[6147] = 8'h0b ;
            rom[6148] = 8'h20 ;
            rom[6149] = 8'hfc ;
            rom[6150] = 8'hf8 ;
            rom[6151] = 8'h0c ;
            rom[6152] = 8'hf4 ;
            rom[6153] = 8'hc7 ;
            rom[6154] = 8'hea ;
            rom[6155] = 8'he2 ;
            rom[6156] = 8'h07 ;
            rom[6157] = 8'h16 ;
            rom[6158] = 8'h1e ;
            rom[6159] = 8'h14 ;
            rom[6160] = 8'h14 ;
            rom[6161] = 8'hf1 ;
            rom[6162] = 8'he4 ;
            rom[6163] = 8'h00 ;
            rom[6164] = 8'hf8 ;
            rom[6165] = 8'h09 ;
            rom[6166] = 8'hfb ;
            rom[6167] = 8'h08 ;
            rom[6168] = 8'hf8 ;
            rom[6169] = 8'hdb ;
            rom[6170] = 8'h29 ;
            rom[6171] = 8'hfa ;
            rom[6172] = 8'he7 ;
            rom[6173] = 8'hf6 ;
            rom[6174] = 8'hec ;
            rom[6175] = 8'hfe ;
            rom[6176] = 8'h0c ;
            rom[6177] = 8'h01 ;
            rom[6178] = 8'h1e ;
            rom[6179] = 8'hd3 ;
            rom[6180] = 8'hec ;
            rom[6181] = 8'hdc ;
            rom[6182] = 8'hed ;
            rom[6183] = 8'h0e ;
            rom[6184] = 8'h06 ;
            rom[6185] = 8'h0d ;
            rom[6186] = 8'hf6 ;
            rom[6187] = 8'heb ;
            rom[6188] = 8'hd6 ;
            rom[6189] = 8'h1d ;
            rom[6190] = 8'hf1 ;
            rom[6191] = 8'hce ;
            rom[6192] = 8'h08 ;
            rom[6193] = 8'hdc ;
            rom[6194] = 8'hea ;
            rom[6195] = 8'hfb ;
            rom[6196] = 8'hf2 ;
            rom[6197] = 8'h0a ;
            rom[6198] = 8'h23 ;
            rom[6199] = 8'h2f ;
            rom[6200] = 8'he0 ;
            rom[6201] = 8'h14 ;
            rom[6202] = 8'h14 ;
            rom[6203] = 8'hed ;
            rom[6204] = 8'hdf ;
            rom[6205] = 8'hb4 ;
            rom[6206] = 8'he7 ;
            rom[6207] = 8'hf0 ;
            rom[6208] = 8'hf2 ;
            rom[6209] = 8'hf4 ;
            rom[6210] = 8'hef ;
            rom[6211] = 8'h0c ;
            rom[6212] = 8'he6 ;
            rom[6213] = 8'hf2 ;
            rom[6214] = 8'h11 ;
            rom[6215] = 8'h14 ;
            rom[6216] = 8'h0f ;
            rom[6217] = 8'h9e ;
            rom[6218] = 8'h06 ;
            rom[6219] = 8'h12 ;
            rom[6220] = 8'hfd ;
            rom[6221] = 8'h03 ;
            rom[6222] = 8'he7 ;
            rom[6223] = 8'hf9 ;
            rom[6224] = 8'hfd ;
            rom[6225] = 8'hd1 ;
            rom[6226] = 8'h05 ;
            rom[6227] = 8'h01 ;
            rom[6228] = 8'h06 ;
            rom[6229] = 8'h0e ;
            rom[6230] = 8'hf0 ;
            rom[6231] = 8'h29 ;
            rom[6232] = 8'h10 ;
            rom[6233] = 8'h37 ;
            rom[6234] = 8'h0b ;
            rom[6235] = 8'hfd ;
            rom[6236] = 8'hf5 ;
            rom[6237] = 8'hf5 ;
            rom[6238] = 8'hf5 ;
            rom[6239] = 8'hf7 ;
            rom[6240] = 8'hed ;
            rom[6241] = 8'h08 ;
            rom[6242] = 8'hfd ;
            rom[6243] = 8'he6 ;
            rom[6244] = 8'hdb ;
            rom[6245] = 8'hf6 ;
            rom[6246] = 8'h19 ;
            rom[6247] = 8'hf2 ;
            rom[6248] = 8'h17 ;
            rom[6249] = 8'hdf ;
            rom[6250] = 8'hea ;
            rom[6251] = 8'hf9 ;
            rom[6252] = 8'h11 ;
            rom[6253] = 8'h04 ;
            rom[6254] = 8'hd9 ;
            rom[6255] = 8'h0c ;
            rom[6256] = 8'h14 ;
            rom[6257] = 8'hf5 ;
            rom[6258] = 8'h12 ;
            rom[6259] = 8'h0f ;
            rom[6260] = 8'hdb ;
            rom[6261] = 8'hf2 ;
            rom[6262] = 8'h15 ;
            rom[6263] = 8'hf9 ;
            rom[6264] = 8'h07 ;
            rom[6265] = 8'h0e ;
            rom[6266] = 8'h05 ;
            rom[6267] = 8'h11 ;
            rom[6268] = 8'h03 ;
            rom[6269] = 8'hff ;
            rom[6270] = 8'h08 ;
            rom[6271] = 8'h24 ;
            rom[6272] = 8'hda ;
            rom[6273] = 8'h9a ;
            rom[6274] = 8'h02 ;
            rom[6275] = 8'hf7 ;
            rom[6276] = 8'he6 ;
            rom[6277] = 8'h22 ;
            rom[6278] = 8'h1c ;
            rom[6279] = 8'h0c ;
            rom[6280] = 8'hf9 ;
            rom[6281] = 8'hb5 ;
            rom[6282] = 8'h23 ;
            rom[6283] = 8'he7 ;
            rom[6284] = 8'h04 ;
            rom[6285] = 8'hd6 ;
            rom[6286] = 8'hf8 ;
            rom[6287] = 8'he1 ;
            rom[6288] = 8'heb ;
            rom[6289] = 8'h0b ;
            rom[6290] = 8'h04 ;
            rom[6291] = 8'h1c ;
            rom[6292] = 8'h06 ;
            rom[6293] = 8'he2 ;
            rom[6294] = 8'h0a ;
            rom[6295] = 8'h10 ;
            rom[6296] = 8'h0b ;
            rom[6297] = 8'hf0 ;
            rom[6298] = 8'h03 ;
            rom[6299] = 8'hf2 ;
            rom[6300] = 8'hd0 ;
            rom[6301] = 8'hfd ;
            rom[6302] = 8'hf6 ;
            rom[6303] = 8'h10 ;
            rom[6304] = 8'h0c ;
            rom[6305] = 8'h14 ;
            rom[6306] = 8'h07 ;
            rom[6307] = 8'he0 ;
            rom[6308] = 8'h13 ;
            rom[6309] = 8'heb ;
            rom[6310] = 8'h14 ;
            rom[6311] = 8'hff ;
            rom[6312] = 8'hfc ;
            rom[6313] = 8'heb ;
            rom[6314] = 8'hf9 ;
            rom[6315] = 8'h11 ;
            rom[6316] = 8'hd9 ;
            rom[6317] = 8'h12 ;
            rom[6318] = 8'hdf ;
            rom[6319] = 8'hdc ;
            rom[6320] = 8'hd8 ;
            rom[6321] = 8'h0f ;
            rom[6322] = 8'he8 ;
            rom[6323] = 8'h04 ;
            rom[6324] = 8'hff ;
            rom[6325] = 8'h02 ;
            rom[6326] = 8'hef ;
            rom[6327] = 8'h17 ;
            rom[6328] = 8'he6 ;
            rom[6329] = 8'he4 ;
            rom[6330] = 8'h24 ;
            rom[6331] = 8'hfb ;
            rom[6332] = 8'hf4 ;
            rom[6333] = 8'he2 ;
            rom[6334] = 8'h04 ;
            rom[6335] = 8'h20 ;
            rom[6336] = 8'hdd ;
            rom[6337] = 8'hfa ;
            rom[6338] = 8'hf5 ;
            rom[6339] = 8'h05 ;
            rom[6340] = 8'h0f ;
            rom[6341] = 8'h2a ;
            rom[6342] = 8'h17 ;
            rom[6343] = 8'hd9 ;
            rom[6344] = 8'h04 ;
            rom[6345] = 8'hd6 ;
            rom[6346] = 8'he4 ;
            rom[6347] = 8'he2 ;
            rom[6348] = 8'he7 ;
            rom[6349] = 8'h0b ;
            rom[6350] = 8'h03 ;
            rom[6351] = 8'hd9 ;
            rom[6352] = 8'hf0 ;
            rom[6353] = 8'hd2 ;
            rom[6354] = 8'h12 ;
            rom[6355] = 8'hc8 ;
            rom[6356] = 8'hf3 ;
            rom[6357] = 8'h06 ;
            rom[6358] = 8'hff ;
            rom[6359] = 8'h1c ;
            rom[6360] = 8'hd0 ;
            rom[6361] = 8'h22 ;
            rom[6362] = 8'hcb ;
            rom[6363] = 8'hdb ;
            rom[6364] = 8'hec ;
            rom[6365] = 8'he0 ;
            rom[6366] = 8'h04 ;
            rom[6367] = 8'hf2 ;
            rom[6368] = 8'he8 ;
            rom[6369] = 8'hfd ;
            rom[6370] = 8'he6 ;
            rom[6371] = 8'h08 ;
            rom[6372] = 8'h16 ;
            rom[6373] = 8'h0f ;
            rom[6374] = 8'h0f ;
            rom[6375] = 8'hce ;
            rom[6376] = 8'hf1 ;
            rom[6377] = 8'hdb ;
            rom[6378] = 8'heb ;
            rom[6379] = 8'h07 ;
            rom[6380] = 8'h02 ;
            rom[6381] = 8'hf9 ;
            rom[6382] = 8'h01 ;
            rom[6383] = 8'hd2 ;
            rom[6384] = 8'h07 ;
            rom[6385] = 8'h0e ;
            rom[6386] = 8'h1d ;
            rom[6387] = 8'hdc ;
            rom[6388] = 8'hfd ;
            rom[6389] = 8'h07 ;
            rom[6390] = 8'hd3 ;
            rom[6391] = 8'hd2 ;
            rom[6392] = 8'h0c ;
            rom[6393] = 8'h02 ;
            rom[6394] = 8'h1c ;
            rom[6395] = 8'h1f ;
            rom[6396] = 8'hd6 ;
            rom[6397] = 8'h07 ;
            rom[6398] = 8'hef ;
            rom[6399] = 8'h23 ;
            rom[6400] = 8'hf2 ;
            rom[6401] = 8'h00 ;
            rom[6402] = 8'hfa ;
            rom[6403] = 8'hd2 ;
            rom[6404] = 8'he8 ;
            rom[6405] = 8'hf9 ;
            rom[6406] = 8'h1d ;
            rom[6407] = 8'hf9 ;
            rom[6408] = 8'hd3 ;
            rom[6409] = 8'hff ;
            rom[6410] = 8'hd0 ;
            rom[6411] = 8'h01 ;
            rom[6412] = 8'he4 ;
            rom[6413] = 8'hf8 ;
            rom[6414] = 8'h13 ;
            rom[6415] = 8'h0f ;
            rom[6416] = 8'h1d ;
            rom[6417] = 8'h00 ;
            rom[6418] = 8'hda ;
            rom[6419] = 8'h00 ;
            rom[6420] = 8'h0f ;
            rom[6421] = 8'h1a ;
            rom[6422] = 8'h00 ;
            rom[6423] = 8'he1 ;
            rom[6424] = 8'hc9 ;
            rom[6425] = 8'h08 ;
            rom[6426] = 8'h00 ;
            rom[6427] = 8'hde ;
            rom[6428] = 8'hf3 ;
            rom[6429] = 8'h10 ;
            rom[6430] = 8'h04 ;
            rom[6431] = 8'hf9 ;
            rom[6432] = 8'he9 ;
            rom[6433] = 8'hea ;
            rom[6434] = 8'hfc ;
            rom[6435] = 8'h11 ;
            rom[6436] = 8'he6 ;
            rom[6437] = 8'hf9 ;
            rom[6438] = 8'h0c ;
            rom[6439] = 8'hd0 ;
            rom[6440] = 8'h09 ;
            rom[6441] = 8'hfd ;
            rom[6442] = 8'h29 ;
            rom[6443] = 8'h11 ;
            rom[6444] = 8'h20 ;
            rom[6445] = 8'hfc ;
            rom[6446] = 8'h08 ;
            rom[6447] = 8'hf4 ;
            rom[6448] = 8'hea ;
            rom[6449] = 8'hd5 ;
            rom[6450] = 8'hfe ;
            rom[6451] = 8'hf9 ;
            rom[6452] = 8'h29 ;
            rom[6453] = 8'h11 ;
            rom[6454] = 8'hfd ;
            rom[6455] = 8'h0e ;
            rom[6456] = 8'hfb ;
            rom[6457] = 8'h05 ;
            rom[6458] = 8'h01 ;
            rom[6459] = 8'h01 ;
            rom[6460] = 8'h0a ;
            rom[6461] = 8'he7 ;
            rom[6462] = 8'h05 ;
            rom[6463] = 8'h02 ;
            rom[6464] = 8'hfd ;
            rom[6465] = 8'h1a ;
            rom[6466] = 8'hf9 ;
            rom[6467] = 8'he9 ;
            rom[6468] = 8'hee ;
            rom[6469] = 8'hf4 ;
            rom[6470] = 8'hc6 ;
            rom[6471] = 8'h2f ;
            rom[6472] = 8'hd1 ;
            rom[6473] = 8'h27 ;
            rom[6474] = 8'hfd ;
            rom[6475] = 8'h06 ;
            rom[6476] = 8'h18 ;
            rom[6477] = 8'he8 ;
            rom[6478] = 8'h2d ;
            rom[6479] = 8'h08 ;
            rom[6480] = 8'hdb ;
            rom[6481] = 8'h09 ;
            rom[6482] = 8'h06 ;
            rom[6483] = 8'h04 ;
            rom[6484] = 8'h22 ;
            rom[6485] = 8'h21 ;
            rom[6486] = 8'h08 ;
            rom[6487] = 8'he9 ;
            rom[6488] = 8'hfa ;
            rom[6489] = 8'h17 ;
            rom[6490] = 8'hf3 ;
            rom[6491] = 8'hf5 ;
            rom[6492] = 8'hf1 ;
            rom[6493] = 8'he5 ;
            rom[6494] = 8'he8 ;
            rom[6495] = 8'h0f ;
            rom[6496] = 8'h01 ;
            rom[6497] = 8'h0e ;
            rom[6498] = 8'he9 ;
            rom[6499] = 8'he0 ;
            rom[6500] = 8'h18 ;
            rom[6501] = 8'hae ;
            rom[6502] = 8'hcd ;
            rom[6503] = 8'h2b ;
            rom[6504] = 8'h09 ;
            rom[6505] = 8'h2d ;
            rom[6506] = 8'he5 ;
            rom[6507] = 8'h1b ;
            rom[6508] = 8'hfe ;
            rom[6509] = 8'hd8 ;
            rom[6510] = 8'hef ;
            rom[6511] = 8'h06 ;
            rom[6512] = 8'hf0 ;
            rom[6513] = 8'h11 ;
            rom[6514] = 8'hed ;
            rom[6515] = 8'h2b ;
            rom[6516] = 8'h0b ;
            rom[6517] = 8'he7 ;
            rom[6518] = 8'h13 ;
            rom[6519] = 8'h03 ;
            rom[6520] = 8'hfb ;
            rom[6521] = 8'h19 ;
            rom[6522] = 8'h00 ;
            rom[6523] = 8'hda ;
            rom[6524] = 8'h23 ;
            rom[6525] = 8'h0c ;
            rom[6526] = 8'hf7 ;
            rom[6527] = 8'h0d ;
            rom[6528] = 8'h09 ;
            rom[6529] = 8'he7 ;
            rom[6530] = 8'hd5 ;
            rom[6531] = 8'he2 ;
            rom[6532] = 8'h02 ;
            rom[6533] = 8'hf5 ;
            rom[6534] = 8'hc7 ;
            rom[6535] = 8'h0c ;
            rom[6536] = 8'h19 ;
            rom[6537] = 8'h04 ;
            rom[6538] = 8'h1a ;
            rom[6539] = 8'hdb ;
            rom[6540] = 8'h10 ;
            rom[6541] = 8'hf3 ;
            rom[6542] = 8'h08 ;
            rom[6543] = 8'hfe ;
            rom[6544] = 8'he6 ;
            rom[6545] = 8'h04 ;
            rom[6546] = 8'h09 ;
            rom[6547] = 8'hef ;
            rom[6548] = 8'h07 ;
            rom[6549] = 8'hda ;
            rom[6550] = 8'hef ;
            rom[6551] = 8'h0b ;
            rom[6552] = 8'h27 ;
            rom[6553] = 8'h06 ;
            rom[6554] = 8'hca ;
            rom[6555] = 8'he0 ;
            rom[6556] = 8'h1a ;
            rom[6557] = 8'h1c ;
            rom[6558] = 8'h00 ;
            rom[6559] = 8'h06 ;
            rom[6560] = 8'h09 ;
            rom[6561] = 8'hea ;
            rom[6562] = 8'h06 ;
            rom[6563] = 8'he6 ;
            rom[6564] = 8'h02 ;
            rom[6565] = 8'h07 ;
            rom[6566] = 8'heb ;
            rom[6567] = 8'h01 ;
            rom[6568] = 8'h15 ;
            rom[6569] = 8'hef ;
            rom[6570] = 8'h15 ;
            rom[6571] = 8'h03 ;
            rom[6572] = 8'h1e ;
            rom[6573] = 8'he4 ;
            rom[6574] = 8'h01 ;
            rom[6575] = 8'hcc ;
            rom[6576] = 8'hf3 ;
            rom[6577] = 8'hf4 ;
            rom[6578] = 8'hdc ;
            rom[6579] = 8'h08 ;
            rom[6580] = 8'h09 ;
            rom[6581] = 8'h1c ;
            rom[6582] = 8'h10 ;
            rom[6583] = 8'hd4 ;
            rom[6584] = 8'hf9 ;
            rom[6585] = 8'hf0 ;
            rom[6586] = 8'h1d ;
            rom[6587] = 8'h0b ;
            rom[6588] = 8'h08 ;
            rom[6589] = 8'hd7 ;
            rom[6590] = 8'h0e ;
            rom[6591] = 8'h0c ;
            rom[6592] = 8'hfd ;
            rom[6593] = 8'h1a ;
            rom[6594] = 8'h13 ;
            rom[6595] = 8'h00 ;
            rom[6596] = 8'h0b ;
            rom[6597] = 8'hfc ;
            rom[6598] = 8'h0c ;
            rom[6599] = 8'hfd ;
            rom[6600] = 8'h06 ;
            rom[6601] = 8'hca ;
            rom[6602] = 8'hd4 ;
            rom[6603] = 8'hda ;
            rom[6604] = 8'he4 ;
            rom[6605] = 8'he1 ;
            rom[6606] = 8'h01 ;
            rom[6607] = 8'hf5 ;
            rom[6608] = 8'h09 ;
            rom[6609] = 8'hdb ;
            rom[6610] = 8'hfd ;
            rom[6611] = 8'hf3 ;
            rom[6612] = 8'hc5 ;
            rom[6613] = 8'h10 ;
            rom[6614] = 8'he3 ;
            rom[6615] = 8'hfb ;
            rom[6616] = 8'h18 ;
            rom[6617] = 8'hff ;
            rom[6618] = 8'h04 ;
            rom[6619] = 8'h1a ;
            rom[6620] = 8'h07 ;
            rom[6621] = 8'hfd ;
            rom[6622] = 8'hf0 ;
            rom[6623] = 8'hee ;
            rom[6624] = 8'hea ;
            rom[6625] = 8'h0c ;
            rom[6626] = 8'hd7 ;
            rom[6627] = 8'h07 ;
            rom[6628] = 8'h0d ;
            rom[6629] = 8'hf8 ;
            rom[6630] = 8'hff ;
            rom[6631] = 8'hff ;
            rom[6632] = 8'hdb ;
            rom[6633] = 8'h1a ;
            rom[6634] = 8'h20 ;
            rom[6635] = 8'hf0 ;
            rom[6636] = 8'h10 ;
            rom[6637] = 8'hf1 ;
            rom[6638] = 8'h02 ;
            rom[6639] = 8'hfd ;
            rom[6640] = 8'heb ;
            rom[6641] = 8'h13 ;
            rom[6642] = 8'h0d ;
            rom[6643] = 8'h04 ;
            rom[6644] = 8'h02 ;
            rom[6645] = 8'hf6 ;
            rom[6646] = 8'h0d ;
            rom[6647] = 8'hf0 ;
            rom[6648] = 8'h16 ;
            rom[6649] = 8'hf6 ;
            rom[6650] = 8'h17 ;
            rom[6651] = 8'hcd ;
            rom[6652] = 8'hc2 ;
            rom[6653] = 8'hea ;
            rom[6654] = 8'hef ;
            rom[6655] = 8'hdd ;
            rom[6656] = 8'heb ;
            rom[6657] = 8'hdc ;
            rom[6658] = 8'hf4 ;
            rom[6659] = 8'h1e ;
            rom[6660] = 8'h07 ;
            rom[6661] = 8'hfe ;
            rom[6662] = 8'hfc ;
            rom[6663] = 8'h0e ;
            rom[6664] = 8'h04 ;
            rom[6665] = 8'h0f ;
            rom[6666] = 8'hfb ;
            rom[6667] = 8'h05 ;
            rom[6668] = 8'hf3 ;
            rom[6669] = 8'hcd ;
            rom[6670] = 8'h04 ;
            rom[6671] = 8'h2b ;
            rom[6672] = 8'h1b ;
            rom[6673] = 8'he7 ;
            rom[6674] = 8'h08 ;
            rom[6675] = 8'hfa ;
            rom[6676] = 8'h1c ;
            rom[6677] = 8'hde ;
            rom[6678] = 8'hf1 ;
            rom[6679] = 8'hf5 ;
            rom[6680] = 8'heb ;
            rom[6681] = 8'hf0 ;
            rom[6682] = 8'hff ;
            rom[6683] = 8'he5 ;
            rom[6684] = 8'h16 ;
            rom[6685] = 8'h0e ;
            rom[6686] = 8'heb ;
            rom[6687] = 8'hd4 ;
            rom[6688] = 8'hf5 ;
            rom[6689] = 8'h05 ;
            rom[6690] = 8'hee ;
            rom[6691] = 8'hfe ;
            rom[6692] = 8'h03 ;
            rom[6693] = 8'h12 ;
            rom[6694] = 8'hff ;
            rom[6695] = 8'h12 ;
            rom[6696] = 8'he2 ;
            rom[6697] = 8'h07 ;
            rom[6698] = 8'h21 ;
            rom[6699] = 8'hf4 ;
            rom[6700] = 8'hf9 ;
            rom[6701] = 8'h14 ;
            rom[6702] = 8'hec ;
            rom[6703] = 8'hf3 ;
            rom[6704] = 8'hf3 ;
            rom[6705] = 8'h2c ;
            rom[6706] = 8'hf5 ;
            rom[6707] = 8'h03 ;
            rom[6708] = 8'hf9 ;
            rom[6709] = 8'he9 ;
            rom[6710] = 8'he6 ;
            rom[6711] = 8'hfc ;
            rom[6712] = 8'h1b ;
            rom[6713] = 8'h36 ;
            rom[6714] = 8'he9 ;
            rom[6715] = 8'hfb ;
            rom[6716] = 8'h23 ;
            rom[6717] = 8'h0d ;
            rom[6718] = 8'hf1 ;
            rom[6719] = 8'hef ;
            rom[6720] = 8'h0c ;
            rom[6721] = 8'hfb ;
            rom[6722] = 8'h0f ;
            rom[6723] = 8'he9 ;
            rom[6724] = 8'hdc ;
            rom[6725] = 8'hc9 ;
            rom[6726] = 8'h11 ;
            rom[6727] = 8'hf5 ;
            rom[6728] = 8'hed ;
            rom[6729] = 8'hde ;
            rom[6730] = 8'hfb ;
            rom[6731] = 8'hf3 ;
            rom[6732] = 8'hdc ;
            rom[6733] = 8'hfb ;
            rom[6734] = 8'hf5 ;
            rom[6735] = 8'h1a ;
            rom[6736] = 8'h14 ;
            rom[6737] = 8'hf0 ;
            rom[6738] = 8'hfd ;
            rom[6739] = 8'hf4 ;
            rom[6740] = 8'hf9 ;
            rom[6741] = 8'hd1 ;
            rom[6742] = 8'hf6 ;
            rom[6743] = 8'heb ;
            rom[6744] = 8'h1c ;
            rom[6745] = 8'hef ;
            rom[6746] = 8'h17 ;
            rom[6747] = 8'h08 ;
            rom[6748] = 8'hef ;
            rom[6749] = 8'he6 ;
            rom[6750] = 8'hcd ;
            rom[6751] = 8'h15 ;
            rom[6752] = 8'hf9 ;
            rom[6753] = 8'h00 ;
            rom[6754] = 8'hd7 ;
            rom[6755] = 8'hf1 ;
            rom[6756] = 8'h1a ;
            rom[6757] = 8'he3 ;
            rom[6758] = 8'h0d ;
            rom[6759] = 8'h18 ;
            rom[6760] = 8'hcc ;
            rom[6761] = 8'hfa ;
            rom[6762] = 8'hf1 ;
            rom[6763] = 8'h09 ;
            rom[6764] = 8'hff ;
            rom[6765] = 8'he0 ;
            rom[6766] = 8'hfc ;
            rom[6767] = 8'h07 ;
            rom[6768] = 8'h0d ;
            rom[6769] = 8'hfa ;
            rom[6770] = 8'h26 ;
            rom[6771] = 8'hf5 ;
            rom[6772] = 8'he3 ;
            rom[6773] = 8'h07 ;
            rom[6774] = 8'h0f ;
            rom[6775] = 8'hde ;
            rom[6776] = 8'hef ;
            rom[6777] = 8'hfa ;
            rom[6778] = 8'h0b ;
            rom[6779] = 8'h11 ;
            rom[6780] = 8'hdc ;
            rom[6781] = 8'he6 ;
            rom[6782] = 8'h0b ;
            rom[6783] = 8'hfd ;
            rom[6784] = 8'hce ;
            rom[6785] = 8'h0e ;
            rom[6786] = 8'hd6 ;
            rom[6787] = 8'h1c ;
            rom[6788] = 8'h0f ;
            rom[6789] = 8'h02 ;
            rom[6790] = 8'hed ;
            rom[6791] = 8'hef ;
            rom[6792] = 8'h0b ;
            rom[6793] = 8'hc7 ;
            rom[6794] = 8'hed ;
            rom[6795] = 8'hf1 ;
            rom[6796] = 8'hd0 ;
            rom[6797] = 8'h09 ;
            rom[6798] = 8'h2e ;
            rom[6799] = 8'hef ;
            rom[6800] = 8'h0a ;
            rom[6801] = 8'h00 ;
            rom[6802] = 8'he5 ;
            rom[6803] = 8'hee ;
            rom[6804] = 8'hf1 ;
            rom[6805] = 8'he9 ;
            rom[6806] = 8'hf4 ;
            rom[6807] = 8'h1e ;
            rom[6808] = 8'h0a ;
            rom[6809] = 8'hf0 ;
            rom[6810] = 8'h25 ;
            rom[6811] = 8'h12 ;
            rom[6812] = 8'he2 ;
            rom[6813] = 8'h1d ;
            rom[6814] = 8'hea ;
            rom[6815] = 8'hfc ;
            rom[6816] = 8'h32 ;
            rom[6817] = 8'h14 ;
            rom[6818] = 8'h03 ;
            rom[6819] = 8'hc9 ;
            rom[6820] = 8'hdd ;
            rom[6821] = 8'hf8 ;
            rom[6822] = 8'h1c ;
            rom[6823] = 8'h15 ;
            rom[6824] = 8'h15 ;
            rom[6825] = 8'he7 ;
            rom[6826] = 8'h09 ;
            rom[6827] = 8'h15 ;
            rom[6828] = 8'h14 ;
            rom[6829] = 8'h27 ;
            rom[6830] = 8'hf5 ;
            rom[6831] = 8'h07 ;
            rom[6832] = 8'hcf ;
            rom[6833] = 8'h22 ;
            rom[6834] = 8'h14 ;
            rom[6835] = 8'h01 ;
            rom[6836] = 8'h11 ;
            rom[6837] = 8'h0f ;
            rom[6838] = 8'he9 ;
            rom[6839] = 8'h2b ;
            rom[6840] = 8'h22 ;
            rom[6841] = 8'hfb ;
            rom[6842] = 8'hf6 ;
            rom[6843] = 8'hf3 ;
            rom[6844] = 8'h02 ;
            rom[6845] = 8'h0b ;
            rom[6846] = 8'h01 ;
            rom[6847] = 8'hf0 ;
            rom[6848] = 8'h27 ;
            rom[6849] = 8'hf7 ;
            rom[6850] = 8'hf3 ;
            rom[6851] = 8'he0 ;
            rom[6852] = 8'h29 ;
            rom[6853] = 8'h23 ;
            rom[6854] = 8'hf8 ;
            rom[6855] = 8'hf5 ;
            rom[6856] = 8'h08 ;
            rom[6857] = 8'hcc ;
            rom[6858] = 8'hf0 ;
            rom[6859] = 8'hed ;
            rom[6860] = 8'h18 ;
            rom[6861] = 8'h2b ;
            rom[6862] = 8'hed ;
            rom[6863] = 8'h1d ;
            rom[6864] = 8'he8 ;
            rom[6865] = 8'hf8 ;
            rom[6866] = 8'h1e ;
            rom[6867] = 8'h04 ;
            rom[6868] = 8'h12 ;
            rom[6869] = 8'he3 ;
            rom[6870] = 8'h0f ;
            rom[6871] = 8'h0b ;
            rom[6872] = 8'hef ;
            rom[6873] = 8'h2f ;
            rom[6874] = 8'hf8 ;
            rom[6875] = 8'hea ;
            rom[6876] = 8'hfb ;
            rom[6877] = 8'h08 ;
            rom[6878] = 8'hf5 ;
            rom[6879] = 8'he7 ;
            rom[6880] = 8'h00 ;
            rom[6881] = 8'h09 ;
            rom[6882] = 8'h07 ;
            rom[6883] = 8'h14 ;
            rom[6884] = 8'hcf ;
            rom[6885] = 8'h0e ;
            rom[6886] = 8'h11 ;
            rom[6887] = 8'hd8 ;
            rom[6888] = 8'hed ;
            rom[6889] = 8'hd3 ;
            rom[6890] = 8'h07 ;
            rom[6891] = 8'h2c ;
            rom[6892] = 8'hf1 ;
            rom[6893] = 8'hea ;
            rom[6894] = 8'hee ;
            rom[6895] = 8'h0d ;
            rom[6896] = 8'hf0 ;
            rom[6897] = 8'hf9 ;
            rom[6898] = 8'h14 ;
            rom[6899] = 8'h22 ;
            rom[6900] = 8'h21 ;
            rom[6901] = 8'hee ;
            rom[6902] = 8'hea ;
            rom[6903] = 8'hfe ;
            rom[6904] = 8'he9 ;
            rom[6905] = 8'hf5 ;
            rom[6906] = 8'hf2 ;
            rom[6907] = 8'hf2 ;
            rom[6908] = 8'hf9 ;
            rom[6909] = 8'h07 ;
            rom[6910] = 8'hd7 ;
            rom[6911] = 8'h0a ;
            rom[6912] = 8'hd4 ;
            rom[6913] = 8'hd9 ;
            rom[6914] = 8'h07 ;
            rom[6915] = 8'he9 ;
            rom[6916] = 8'h07 ;
            rom[6917] = 8'h14 ;
            rom[6918] = 8'hd9 ;
            rom[6919] = 8'h05 ;
            rom[6920] = 8'hed ;
            rom[6921] = 8'hed ;
            rom[6922] = 8'h06 ;
            rom[6923] = 8'hdd ;
            rom[6924] = 8'hf3 ;
            rom[6925] = 8'h0f ;
            rom[6926] = 8'h1e ;
            rom[6927] = 8'hf5 ;
            rom[6928] = 8'h03 ;
            rom[6929] = 8'h10 ;
            rom[6930] = 8'he9 ;
            rom[6931] = 8'hfd ;
            rom[6932] = 8'hf3 ;
            rom[6933] = 8'hf4 ;
            rom[6934] = 8'h30 ;
            rom[6935] = 8'hdc ;
            rom[6936] = 8'hc2 ;
            rom[6937] = 8'hf7 ;
            rom[6938] = 8'hf0 ;
            rom[6939] = 8'hf4 ;
            rom[6940] = 8'h08 ;
            rom[6941] = 8'h09 ;
            rom[6942] = 8'hf8 ;
            rom[6943] = 8'h12 ;
            rom[6944] = 8'he4 ;
            rom[6945] = 8'hfe ;
            rom[6946] = 8'hf1 ;
            rom[6947] = 8'h05 ;
            rom[6948] = 8'he1 ;
            rom[6949] = 8'hab ;
            rom[6950] = 8'hf7 ;
            rom[6951] = 8'h08 ;
            rom[6952] = 8'h0f ;
            rom[6953] = 8'hfa ;
            rom[6954] = 8'h16 ;
            rom[6955] = 8'hfd ;
            rom[6956] = 8'he0 ;
            rom[6957] = 8'he0 ;
            rom[6958] = 8'hf6 ;
            rom[6959] = 8'h0e ;
            rom[6960] = 8'hf1 ;
            rom[6961] = 8'hd0 ;
            rom[6962] = 8'h0e ;
            rom[6963] = 8'hec ;
            rom[6964] = 8'hfd ;
            rom[6965] = 8'h0d ;
            rom[6966] = 8'h16 ;
            rom[6967] = 8'h11 ;
            rom[6968] = 8'he3 ;
            rom[6969] = 8'h04 ;
            rom[6970] = 8'h2f ;
            rom[6971] = 8'hd8 ;
            rom[6972] = 8'hf5 ;
            rom[6973] = 8'h0d ;
            rom[6974] = 8'h03 ;
            rom[6975] = 8'hf3 ;
            rom[6976] = 8'h1a ;
            rom[6977] = 8'hfe ;
            rom[6978] = 8'h14 ;
            rom[6979] = 8'h1b ;
            rom[6980] = 8'h07 ;
            rom[6981] = 8'hf9 ;
            rom[6982] = 8'h0a ;
            rom[6983] = 8'h16 ;
            rom[6984] = 8'h0c ;
            rom[6985] = 8'hdf ;
            rom[6986] = 8'hf9 ;
            rom[6987] = 8'h13 ;
            rom[6988] = 8'h01 ;
            rom[6989] = 8'hec ;
            rom[6990] = 8'h12 ;
            rom[6991] = 8'hfd ;
            rom[6992] = 8'h12 ;
            rom[6993] = 8'hea ;
            rom[6994] = 8'h05 ;
            rom[6995] = 8'hd8 ;
            rom[6996] = 8'h08 ;
            rom[6997] = 8'hf2 ;
            rom[6998] = 8'h0e ;
            rom[6999] = 8'h0f ;
            rom[7000] = 8'hed ;
            rom[7001] = 8'h11 ;
            rom[7002] = 8'hf0 ;
            rom[7003] = 8'he4 ;
            rom[7004] = 8'hdc ;
            rom[7005] = 8'he0 ;
            rom[7006] = 8'hf4 ;
            rom[7007] = 8'hef ;
            rom[7008] = 8'hd5 ;
            rom[7009] = 8'hf4 ;
            rom[7010] = 8'he4 ;
            rom[7011] = 8'heb ;
            rom[7012] = 8'hed ;
            rom[7013] = 8'hd1 ;
            rom[7014] = 8'hf8 ;
            rom[7015] = 8'h09 ;
            rom[7016] = 8'hfe ;
            rom[7017] = 8'h21 ;
            rom[7018] = 8'hfc ;
            rom[7019] = 8'h0b ;
            rom[7020] = 8'h1c ;
            rom[7021] = 8'h09 ;
            rom[7022] = 8'h0e ;
            rom[7023] = 8'he3 ;
            rom[7024] = 8'he3 ;
            rom[7025] = 8'h03 ;
            rom[7026] = 8'h22 ;
            rom[7027] = 8'h1f ;
            rom[7028] = 8'hdb ;
            rom[7029] = 8'h1a ;
            rom[7030] = 8'h0f ;
            rom[7031] = 8'h10 ;
            rom[7032] = 8'h20 ;
            rom[7033] = 8'hf1 ;
            rom[7034] = 8'h27 ;
            rom[7035] = 8'hd1 ;
            rom[7036] = 8'he3 ;
            rom[7037] = 8'hf9 ;
            rom[7038] = 8'hf8 ;
            rom[7039] = 8'hcb ;
            rom[7040] = 8'he3 ;
            rom[7041] = 8'hd7 ;
            rom[7042] = 8'h03 ;
            rom[7043] = 8'h0a ;
            rom[7044] = 8'hfa ;
            rom[7045] = 8'hf8 ;
            rom[7046] = 8'h14 ;
            rom[7047] = 8'hcd ;
            rom[7048] = 8'hef ;
            rom[7049] = 8'h07 ;
            rom[7050] = 8'hec ;
            rom[7051] = 8'h1e ;
            rom[7052] = 8'hef ;
            rom[7053] = 8'hff ;
            rom[7054] = 8'hc7 ;
            rom[7055] = 8'hfc ;
            rom[7056] = 8'hf9 ;
            rom[7057] = 8'h27 ;
            rom[7058] = 8'h18 ;
            rom[7059] = 8'hf4 ;
            rom[7060] = 8'h12 ;
            rom[7061] = 8'h0a ;
            rom[7062] = 8'hde ;
            rom[7063] = 8'hec ;
            rom[7064] = 8'hea ;
            rom[7065] = 8'h12 ;
            rom[7066] = 8'h23 ;
            rom[7067] = 8'hf9 ;
            rom[7068] = 8'hcb ;
            rom[7069] = 8'h04 ;
            rom[7070] = 8'hee ;
            rom[7071] = 8'h02 ;
            rom[7072] = 8'hf2 ;
            rom[7073] = 8'hf3 ;
            rom[7074] = 8'hef ;
            rom[7075] = 8'h15 ;
            rom[7076] = 8'h09 ;
            rom[7077] = 8'h04 ;
            rom[7078] = 8'h0b ;
            rom[7079] = 8'h1b ;
            rom[7080] = 8'h11 ;
            rom[7081] = 8'hfb ;
            rom[7082] = 8'h19 ;
            rom[7083] = 8'hff ;
            rom[7084] = 8'hfd ;
            rom[7085] = 8'hff ;
            rom[7086] = 8'hfd ;
            rom[7087] = 8'hfd ;
            rom[7088] = 8'hd5 ;
            rom[7089] = 8'h00 ;
            rom[7090] = 8'h15 ;
            rom[7091] = 8'hdb ;
            rom[7092] = 8'h12 ;
            rom[7093] = 8'hcc ;
            rom[7094] = 8'hdd ;
            rom[7095] = 8'h1d ;
            rom[7096] = 8'h39 ;
            rom[7097] = 8'h0c ;
            rom[7098] = 8'hfd ;
            rom[7099] = 8'hfe ;
            rom[7100] = 8'h19 ;
            rom[7101] = 8'hf3 ;
            rom[7102] = 8'h05 ;
            rom[7103] = 8'h01 ;
            rom[7104] = 8'hf6 ;
            rom[7105] = 8'he2 ;
            rom[7106] = 8'h12 ;
            rom[7107] = 8'hdb ;
            rom[7108] = 8'hf1 ;
            rom[7109] = 8'he9 ;
            rom[7110] = 8'hd8 ;
            rom[7111] = 8'hed ;
            rom[7112] = 8'he4 ;
            rom[7113] = 8'h0f ;
            rom[7114] = 8'h1b ;
            rom[7115] = 8'he0 ;
            rom[7116] = 8'h0f ;
            rom[7117] = 8'hf2 ;
            rom[7118] = 8'h1d ;
            rom[7119] = 8'h09 ;
            rom[7120] = 8'hd8 ;
            rom[7121] = 8'h22 ;
            rom[7122] = 8'hc9 ;
            rom[7123] = 8'hfb ;
            rom[7124] = 8'h00 ;
            rom[7125] = 8'hed ;
            rom[7126] = 8'hff ;
            rom[7127] = 8'he5 ;
            rom[7128] = 8'h08 ;
            rom[7129] = 8'h1b ;
            rom[7130] = 8'hd7 ;
            rom[7131] = 8'hdb ;
            rom[7132] = 8'hf6 ;
            rom[7133] = 8'h14 ;
            rom[7134] = 8'h1e ;
            rom[7135] = 8'h0d ;
            rom[7136] = 8'hff ;
            rom[7137] = 8'he3 ;
            rom[7138] = 8'h04 ;
            rom[7139] = 8'h11 ;
            rom[7140] = 8'heb ;
            rom[7141] = 8'hd0 ;
            rom[7142] = 8'hd9 ;
            rom[7143] = 8'hce ;
            rom[7144] = 8'hf9 ;
            rom[7145] = 8'h05 ;
            rom[7146] = 8'hdd ;
            rom[7147] = 8'hf3 ;
            rom[7148] = 8'hc9 ;
            rom[7149] = 8'hda ;
            rom[7150] = 8'h1a ;
            rom[7151] = 8'hea ;
            rom[7152] = 8'he6 ;
            rom[7153] = 8'h1c ;
            rom[7154] = 8'h03 ;
            rom[7155] = 8'h1d ;
            rom[7156] = 8'h03 ;
            rom[7157] = 8'hef ;
            rom[7158] = 8'hf4 ;
            rom[7159] = 8'h10 ;
            rom[7160] = 8'he2 ;
            rom[7161] = 8'h1a ;
            rom[7162] = 8'hed ;
            rom[7163] = 8'h0e ;
            rom[7164] = 8'hfc ;
            rom[7165] = 8'hf5 ;
            rom[7166] = 8'hc1 ;
            rom[7167] = 8'h19 ;
            rom[7168] = 8'hf6 ;
            rom[7169] = 8'h03 ;
            rom[7170] = 8'h26 ;
            rom[7171] = 8'hfa ;
            rom[7172] = 8'hee ;
            rom[7173] = 8'hef ;
            rom[7174] = 8'h0b ;
            rom[7175] = 8'hf7 ;
            rom[7176] = 8'h0d ;
            rom[7177] = 8'hdd ;
            rom[7178] = 8'hf6 ;
            rom[7179] = 8'h1f ;
            rom[7180] = 8'hf5 ;
            rom[7181] = 8'hde ;
            rom[7182] = 8'hdf ;
            rom[7183] = 8'h10 ;
            rom[7184] = 8'h00 ;
            rom[7185] = 8'he7 ;
            rom[7186] = 8'h07 ;
            rom[7187] = 8'h1d ;
            rom[7188] = 8'hf7 ;
            rom[7189] = 8'he9 ;
            rom[7190] = 8'h26 ;
            rom[7191] = 8'h1d ;
            rom[7192] = 8'hf6 ;
            rom[7193] = 8'heb ;
            rom[7194] = 8'h07 ;
            rom[7195] = 8'h12 ;
            rom[7196] = 8'hd5 ;
            rom[7197] = 8'h05 ;
            rom[7198] = 8'hd2 ;
            rom[7199] = 8'hdb ;
            rom[7200] = 8'hdd ;
            rom[7201] = 8'hf8 ;
            rom[7202] = 8'hf4 ;
            rom[7203] = 8'hcc ;
            rom[7204] = 8'hf8 ;
            rom[7205] = 8'hfb ;
            rom[7206] = 8'hed ;
            rom[7207] = 8'he4 ;
            rom[7208] = 8'h06 ;
            rom[7209] = 8'heb ;
            rom[7210] = 8'h20 ;
            rom[7211] = 8'h19 ;
            rom[7212] = 8'he6 ;
            rom[7213] = 8'h10 ;
            rom[7214] = 8'hf9 ;
            rom[7215] = 8'hf1 ;
            rom[7216] = 8'hfa ;
            rom[7217] = 8'h17 ;
            rom[7218] = 8'hdc ;
            rom[7219] = 8'h06 ;
            rom[7220] = 8'hfb ;
            rom[7221] = 8'he4 ;
            rom[7222] = 8'heb ;
            rom[7223] = 8'h09 ;
            rom[7224] = 8'hfc ;
            rom[7225] = 8'hf3 ;
            rom[7226] = 8'h01 ;
            rom[7227] = 8'h0a ;
            rom[7228] = 8'h33 ;
            rom[7229] = 8'hed ;
            rom[7230] = 8'h16 ;
            rom[7231] = 8'hdb ;
            rom[7232] = 8'h05 ;
            rom[7233] = 8'h17 ;
            rom[7234] = 8'he1 ;
            rom[7235] = 8'hfa ;
            rom[7236] = 8'he5 ;
            rom[7237] = 8'h12 ;
            rom[7238] = 8'hfb ;
            rom[7239] = 8'hbb ;
            rom[7240] = 8'hfc ;
            rom[7241] = 8'h0f ;
            rom[7242] = 8'hed ;
            rom[7243] = 8'h03 ;
            rom[7244] = 8'hdd ;
            rom[7245] = 8'h18 ;
            rom[7246] = 8'h07 ;
            rom[7247] = 8'hef ;
            rom[7248] = 8'hd7 ;
            rom[7249] = 8'h0f ;
            rom[7250] = 8'hf4 ;
            rom[7251] = 8'hf5 ;
            rom[7252] = 8'hed ;
            rom[7253] = 8'he6 ;
            rom[7254] = 8'hf6 ;
            rom[7255] = 8'hd7 ;
            rom[7256] = 8'hf8 ;
            rom[7257] = 8'hf1 ;
            rom[7258] = 8'h08 ;
            rom[7259] = 8'he6 ;
            rom[7260] = 8'hf8 ;
            rom[7261] = 8'hf0 ;
            rom[7262] = 8'h11 ;
            rom[7263] = 8'hba ;
            rom[7264] = 8'h12 ;
            rom[7265] = 8'h0d ;
            rom[7266] = 8'he0 ;
            rom[7267] = 8'h1c ;
            rom[7268] = 8'h0d ;
            rom[7269] = 8'hee ;
            rom[7270] = 8'he8 ;
            rom[7271] = 8'hf3 ;
            rom[7272] = 8'he1 ;
            rom[7273] = 8'hf1 ;
            rom[7274] = 8'he6 ;
            rom[7275] = 8'h29 ;
            rom[7276] = 8'he5 ;
            rom[7277] = 8'h04 ;
            rom[7278] = 8'he3 ;
            rom[7279] = 8'hfd ;
            rom[7280] = 8'he0 ;
            rom[7281] = 8'h09 ;
            rom[7282] = 8'h05 ;
            rom[7283] = 8'he0 ;
            rom[7284] = 8'h03 ;
            rom[7285] = 8'hf3 ;
            rom[7286] = 8'hbf ;
            rom[7287] = 8'he2 ;
            rom[7288] = 8'hfe ;
            rom[7289] = 8'hce ;
            rom[7290] = 8'hf1 ;
            rom[7291] = 8'h11 ;
            rom[7292] = 8'hf3 ;
            rom[7293] = 8'he1 ;
            rom[7294] = 8'hf5 ;
            rom[7295] = 8'hee ;
            rom[7296] = 8'hfc ;
            rom[7297] = 8'h08 ;
            rom[7298] = 8'hf1 ;
            rom[7299] = 8'h05 ;
            rom[7300] = 8'hfd ;
            rom[7301] = 8'h1f ;
            rom[7302] = 8'hdf ;
            rom[7303] = 8'h1a ;
            rom[7304] = 8'hf4 ;
            rom[7305] = 8'h03 ;
            rom[7306] = 8'hfe ;
            rom[7307] = 8'hdb ;
            rom[7308] = 8'he9 ;
            rom[7309] = 8'hfa ;
            rom[7310] = 8'h18 ;
            rom[7311] = 8'he6 ;
            rom[7312] = 8'h2d ;
            rom[7313] = 8'h10 ;
            rom[7314] = 8'he6 ;
            rom[7315] = 8'h09 ;
            rom[7316] = 8'hfe ;
            rom[7317] = 8'hfb ;
            rom[7318] = 8'hf2 ;
            rom[7319] = 8'hfe ;
            rom[7320] = 8'h04 ;
            rom[7321] = 8'hf9 ;
            rom[7322] = 8'h04 ;
            rom[7323] = 8'hea ;
            rom[7324] = 8'h05 ;
            rom[7325] = 8'h21 ;
            rom[7326] = 8'hf5 ;
            rom[7327] = 8'h09 ;
            rom[7328] = 8'hde ;
            rom[7329] = 8'h16 ;
            rom[7330] = 8'he4 ;
            rom[7331] = 8'h22 ;
            rom[7332] = 8'hfb ;
            rom[7333] = 8'hc4 ;
            rom[7334] = 8'h0b ;
            rom[7335] = 8'hf4 ;
            rom[7336] = 8'h0c ;
            rom[7337] = 8'h02 ;
            rom[7338] = 8'h0d ;
            rom[7339] = 8'hff ;
            rom[7340] = 8'h15 ;
            rom[7341] = 8'hce ;
            rom[7342] = 8'h06 ;
            rom[7343] = 8'hdf ;
            rom[7344] = 8'hef ;
            rom[7345] = 8'hdc ;
            rom[7346] = 8'h01 ;
            rom[7347] = 8'h08 ;
            rom[7348] = 8'h12 ;
            rom[7349] = 8'hf3 ;
            rom[7350] = 8'he8 ;
            rom[7351] = 8'h10 ;
            rom[7352] = 8'h1c ;
            rom[7353] = 8'h04 ;
            rom[7354] = 8'h00 ;
            rom[7355] = 8'hf6 ;
            rom[7356] = 8'hf9 ;
            rom[7357] = 8'hdf ;
            rom[7358] = 8'h2a ;
            rom[7359] = 8'h16 ;
            rom[7360] = 8'hfc ;
            rom[7361] = 8'h20 ;
            rom[7362] = 8'h16 ;
            rom[7363] = 8'hef ;
            rom[7364] = 8'hf0 ;
            rom[7365] = 8'heb ;
            rom[7366] = 8'h0a ;
            rom[7367] = 8'h1f ;
            rom[7368] = 8'h12 ;
            rom[7369] = 8'h00 ;
            rom[7370] = 8'h19 ;
            rom[7371] = 8'h07 ;
            rom[7372] = 8'h0e ;
            rom[7373] = 8'h06 ;
            rom[7374] = 8'h22 ;
            rom[7375] = 8'h11 ;
            rom[7376] = 8'h11 ;
            rom[7377] = 8'h06 ;
            rom[7378] = 8'hfc ;
            rom[7379] = 8'he6 ;
            rom[7380] = 8'hfd ;
            rom[7381] = 8'h35 ;
            rom[7382] = 8'hf1 ;
            rom[7383] = 8'h14 ;
            rom[7384] = 8'he7 ;
            rom[7385] = 8'h27 ;
            rom[7386] = 8'he3 ;
            rom[7387] = 8'hfd ;
            rom[7388] = 8'hea ;
            rom[7389] = 8'h02 ;
            rom[7390] = 8'hd4 ;
            rom[7391] = 8'h13 ;
            rom[7392] = 8'hf6 ;
            rom[7393] = 8'h05 ;
            rom[7394] = 8'h08 ;
            rom[7395] = 8'hde ;
            rom[7396] = 8'heb ;
            rom[7397] = 8'hca ;
            rom[7398] = 8'h04 ;
            rom[7399] = 8'h04 ;
            rom[7400] = 8'hf2 ;
            rom[7401] = 8'h06 ;
            rom[7402] = 8'he0 ;
            rom[7403] = 8'h20 ;
            rom[7404] = 8'h09 ;
            rom[7405] = 8'hbc ;
            rom[7406] = 8'h11 ;
            rom[7407] = 8'h07 ;
            rom[7408] = 8'hc6 ;
            rom[7409] = 8'h06 ;
            rom[7410] = 8'hd3 ;
            rom[7411] = 8'h2f ;
            rom[7412] = 8'h22 ;
            rom[7413] = 8'hdf ;
            rom[7414] = 8'h30 ;
            rom[7415] = 8'h22 ;
            rom[7416] = 8'h18 ;
            rom[7417] = 8'h04 ;
            rom[7418] = 8'h13 ;
            rom[7419] = 8'hd0 ;
            rom[7420] = 8'h03 ;
            rom[7421] = 8'h07 ;
            rom[7422] = 8'h0b ;
            rom[7423] = 8'h1f ;
            rom[7424] = 8'h27 ;
            rom[7425] = 8'h08 ;
            rom[7426] = 8'hf5 ;
            rom[7427] = 8'h14 ;
            rom[7428] = 8'hff ;
            rom[7429] = 8'hff ;
            rom[7430] = 8'hf9 ;
            rom[7431] = 8'hed ;
            rom[7432] = 8'he5 ;
            rom[7433] = 8'h20 ;
            rom[7434] = 8'h27 ;
            rom[7435] = 8'hce ;
            rom[7436] = 8'hcb ;
            rom[7437] = 8'hf9 ;
            rom[7438] = 8'h26 ;
            rom[7439] = 8'hbe ;
            rom[7440] = 8'hd8 ;
            rom[7441] = 8'hf3 ;
            rom[7442] = 8'hce ;
            rom[7443] = 8'h01 ;
            rom[7444] = 8'hfe ;
            rom[7445] = 8'hcd ;
            rom[7446] = 8'h17 ;
            rom[7447] = 8'h06 ;
            rom[7448] = 8'h02 ;
            rom[7449] = 8'h07 ;
            rom[7450] = 8'hf7 ;
            rom[7451] = 8'hda ;
            rom[7452] = 8'h1c ;
            rom[7453] = 8'h1d ;
            rom[7454] = 8'h02 ;
            rom[7455] = 8'h12 ;
            rom[7456] = 8'he6 ;
            rom[7457] = 8'h19 ;
            rom[7458] = 8'h1b ;
            rom[7459] = 8'hdf ;
            rom[7460] = 8'h29 ;
            rom[7461] = 8'hfc ;
            rom[7462] = 8'he7 ;
            rom[7463] = 8'h0f ;
            rom[7464] = 8'hf2 ;
            rom[7465] = 8'hff ;
            rom[7466] = 8'hf7 ;
            rom[7467] = 8'hfc ;
            rom[7468] = 8'hfa ;
            rom[7469] = 8'hfb ;
            rom[7470] = 8'hfc ;
            rom[7471] = 8'hed ;
            rom[7472] = 8'hfd ;
            rom[7473] = 8'h0e ;
            rom[7474] = 8'hcb ;
            rom[7475] = 8'hef ;
            rom[7476] = 8'h02 ;
            rom[7477] = 8'h02 ;
            rom[7478] = 8'hea ;
            rom[7479] = 8'he7 ;
            rom[7480] = 8'h0d ;
            rom[7481] = 8'h05 ;
            rom[7482] = 8'h07 ;
            rom[7483] = 8'hda ;
            rom[7484] = 8'h00 ;
            rom[7485] = 8'he1 ;
            rom[7486] = 8'h0a ;
            rom[7487] = 8'h02 ;
            rom[7488] = 8'h05 ;
            rom[7489] = 8'hff ;
            rom[7490] = 8'h28 ;
            rom[7491] = 8'hbf ;
            rom[7492] = 8'h12 ;
            rom[7493] = 8'hfc ;
            rom[7494] = 8'he6 ;
            rom[7495] = 8'he2 ;
            rom[7496] = 8'h18 ;
            rom[7497] = 8'hfd ;
            rom[7498] = 8'hdd ;
            rom[7499] = 8'hce ;
            rom[7500] = 8'he1 ;
            rom[7501] = 8'he2 ;
            rom[7502] = 8'he9 ;
            rom[7503] = 8'h13 ;
            rom[7504] = 8'h1a ;
            rom[7505] = 8'hf3 ;
            rom[7506] = 8'h1b ;
            rom[7507] = 8'hcd ;
            rom[7508] = 8'hdb ;
            rom[7509] = 8'h0e ;
            rom[7510] = 8'hd3 ;
            rom[7511] = 8'h06 ;
            rom[7512] = 8'h0b ;
            rom[7513] = 8'hf1 ;
            rom[7514] = 8'hfe ;
            rom[7515] = 8'hf9 ;
            rom[7516] = 8'hd7 ;
            rom[7517] = 8'h02 ;
            rom[7518] = 8'h08 ;
            rom[7519] = 8'hd8 ;
            rom[7520] = 8'he6 ;
            rom[7521] = 8'heb ;
            rom[7522] = 8'h06 ;
            rom[7523] = 8'h02 ;
            rom[7524] = 8'h08 ;
            rom[7525] = 8'h1d ;
            rom[7526] = 8'h0a ;
            rom[7527] = 8'hf9 ;
            rom[7528] = 8'hc9 ;
            rom[7529] = 8'hf4 ;
            rom[7530] = 8'h22 ;
            rom[7531] = 8'hef ;
            rom[7532] = 8'h13 ;
            rom[7533] = 8'hfd ;
            rom[7534] = 8'h05 ;
            rom[7535] = 8'h01 ;
            rom[7536] = 8'hdf ;
            rom[7537] = 8'hfd ;
            rom[7538] = 8'hf2 ;
            rom[7539] = 8'hf9 ;
            rom[7540] = 8'h00 ;
            rom[7541] = 8'h14 ;
            rom[7542] = 8'he1 ;
            rom[7543] = 8'hff ;
            rom[7544] = 8'he3 ;
            rom[7545] = 8'hdb ;
            rom[7546] = 8'hf4 ;
            rom[7547] = 8'h1b ;
            rom[7548] = 8'hcd ;
            rom[7549] = 8'h0b ;
            rom[7550] = 8'h0d ;
            rom[7551] = 8'hf2 ;
            rom[7552] = 8'hef ;
            rom[7553] = 8'hfc ;
            rom[7554] = 8'hf3 ;
            rom[7555] = 8'h0a ;
            rom[7556] = 8'h1b ;
            rom[7557] = 8'hdb ;
            rom[7558] = 8'hf4 ;
            rom[7559] = 8'hf1 ;
            rom[7560] = 8'he5 ;
            rom[7561] = 8'h11 ;
            rom[7562] = 8'hfe ;
            rom[7563] = 8'hdc ;
            rom[7564] = 8'hec ;
            rom[7565] = 8'h0e ;
            rom[7566] = 8'hee ;
            rom[7567] = 8'h15 ;
            rom[7568] = 8'hfa ;
            rom[7569] = 8'h17 ;
            rom[7570] = 8'he7 ;
            rom[7571] = 8'hd7 ;
            rom[7572] = 8'h1a ;
            rom[7573] = 8'h11 ;
            rom[7574] = 8'h03 ;
            rom[7575] = 8'hfb ;
            rom[7576] = 8'hd3 ;
            rom[7577] = 8'h12 ;
            rom[7578] = 8'h01 ;
            rom[7579] = 8'h18 ;
            rom[7580] = 8'h04 ;
            rom[7581] = 8'h04 ;
            rom[7582] = 8'hf6 ;
            rom[7583] = 8'hf2 ;
            rom[7584] = 8'h22 ;
            rom[7585] = 8'he2 ;
            rom[7586] = 8'hc7 ;
            rom[7587] = 8'he3 ;
            rom[7588] = 8'hde ;
            rom[7589] = 8'hd1 ;
            rom[7590] = 8'h12 ;
            rom[7591] = 8'hff ;
            rom[7592] = 8'h16 ;
            rom[7593] = 8'hf8 ;
            rom[7594] = 8'hf3 ;
            rom[7595] = 8'h04 ;
            rom[7596] = 8'h01 ;
            rom[7597] = 8'hd2 ;
            rom[7598] = 8'h01 ;
            rom[7599] = 8'h17 ;
            rom[7600] = 8'hfc ;
            rom[7601] = 8'h03 ;
            rom[7602] = 8'h26 ;
            rom[7603] = 8'hf5 ;
            rom[7604] = 8'h15 ;
            rom[7605] = 8'hf8 ;
            rom[7606] = 8'he8 ;
            rom[7607] = 8'hf2 ;
            rom[7608] = 8'h0c ;
            rom[7609] = 8'hf8 ;
            rom[7610] = 8'h14 ;
            rom[7611] = 8'hfc ;
            rom[7612] = 8'hed ;
            rom[7613] = 8'h09 ;
            rom[7614] = 8'hf8 ;
            rom[7615] = 8'hf2 ;
            rom[7616] = 8'h18 ;
            rom[7617] = 8'h23 ;
            rom[7618] = 8'h06 ;
            rom[7619] = 8'hc6 ;
            rom[7620] = 8'h04 ;
            rom[7621] = 8'he2 ;
            rom[7622] = 8'hf3 ;
            rom[7623] = 8'h00 ;
            rom[7624] = 8'h27 ;
            rom[7625] = 8'hf3 ;
            rom[7626] = 8'h15 ;
            rom[7627] = 8'hf8 ;
            rom[7628] = 8'h00 ;
            rom[7629] = 8'hf9 ;
            rom[7630] = 8'hf4 ;
            rom[7631] = 8'h11 ;
            rom[7632] = 8'hb4 ;
            rom[7633] = 8'h0b ;
            rom[7634] = 8'hf3 ;
            rom[7635] = 8'h0e ;
            rom[7636] = 8'h11 ;
            rom[7637] = 8'h22 ;
            rom[7638] = 8'h16 ;
            rom[7639] = 8'heb ;
            rom[7640] = 8'h0a ;
            rom[7641] = 8'h14 ;
            rom[7642] = 8'h05 ;
            rom[7643] = 8'h08 ;
            rom[7644] = 8'hee ;
            rom[7645] = 8'h19 ;
            rom[7646] = 8'h02 ;
            rom[7647] = 8'h25 ;
            rom[7648] = 8'he6 ;
            rom[7649] = 8'hef ;
            rom[7650] = 8'hf4 ;
            rom[7651] = 8'hea ;
            rom[7652] = 8'h1c ;
            rom[7653] = 8'hb4 ;
            rom[7654] = 8'hea ;
            rom[7655] = 8'h04 ;
            rom[7656] = 8'hd4 ;
            rom[7657] = 8'h31 ;
            rom[7658] = 8'he9 ;
            rom[7659] = 8'hf0 ;
            rom[7660] = 8'ha1 ;
            rom[7661] = 8'hde ;
            rom[7662] = 8'hcc ;
            rom[7663] = 8'h20 ;
            rom[7664] = 8'hf7 ;
            rom[7665] = 8'h02 ;
            rom[7666] = 8'h01 ;
            rom[7667] = 8'h2b ;
            rom[7668] = 8'h12 ;
            rom[7669] = 8'h04 ;
            rom[7670] = 8'hf9 ;
            rom[7671] = 8'h24 ;
            rom[7672] = 8'hfe ;
            rom[7673] = 8'hf8 ;
            rom[7674] = 8'hdf ;
            rom[7675] = 8'h04 ;
            rom[7676] = 8'h04 ;
            rom[7677] = 8'h0a ;
            rom[7678] = 8'hc8 ;
            rom[7679] = 8'he1 ;
            rom[7680] = 8'hd2 ;
            rom[7681] = 8'hdf ;
            rom[7682] = 8'hfa ;
            rom[7683] = 8'h13 ;
            rom[7684] = 8'h03 ;
            rom[7685] = 8'hfe ;
            rom[7686] = 8'he6 ;
            rom[7687] = 8'hfa ;
            rom[7688] = 8'hd9 ;
            rom[7689] = 8'h1f ;
            rom[7690] = 8'h1a ;
            rom[7691] = 8'hfa ;
            rom[7692] = 8'hef ;
            rom[7693] = 8'h09 ;
            rom[7694] = 8'hfd ;
            rom[7695] = 8'h0f ;
            rom[7696] = 8'h0f ;
            rom[7697] = 8'h17 ;
            rom[7698] = 8'hd6 ;
            rom[7699] = 8'hea ;
            rom[7700] = 8'h10 ;
            rom[7701] = 8'h08 ;
            rom[7702] = 8'hd8 ;
            rom[7703] = 8'h22 ;
            rom[7704] = 8'h01 ;
            rom[7705] = 8'h1d ;
            rom[7706] = 8'hff ;
            rom[7707] = 8'h0b ;
            rom[7708] = 8'he6 ;
            rom[7709] = 8'h1c ;
            rom[7710] = 8'h11 ;
            rom[7711] = 8'h07 ;
            rom[7712] = 8'he6 ;
            rom[7713] = 8'h15 ;
            rom[7714] = 8'h12 ;
            rom[7715] = 8'h00 ;
            rom[7716] = 8'hf9 ;
            rom[7717] = 8'h04 ;
            rom[7718] = 8'h01 ;
            rom[7719] = 8'h0d ;
            rom[7720] = 8'hef ;
            rom[7721] = 8'hf0 ;
            rom[7722] = 8'hd7 ;
            rom[7723] = 8'hf7 ;
            rom[7724] = 8'hf9 ;
            rom[7725] = 8'hdf ;
            rom[7726] = 8'hff ;
            rom[7727] = 8'he7 ;
            rom[7728] = 8'hd1 ;
            rom[7729] = 8'hd7 ;
            rom[7730] = 8'hfc ;
            rom[7731] = 8'hde ;
            rom[7732] = 8'h1c ;
            rom[7733] = 8'he0 ;
            rom[7734] = 8'h1d ;
            rom[7735] = 8'hf6 ;
            rom[7736] = 8'h1e ;
            rom[7737] = 8'hf6 ;
            rom[7738] = 8'h06 ;
            rom[7739] = 8'hc9 ;
            rom[7740] = 8'h17 ;
            rom[7741] = 8'he4 ;
            rom[7742] = 8'hfb ;
            rom[7743] = 8'h07 ;
            rom[7744] = 8'h21 ;
            rom[7745] = 8'h04 ;
            rom[7746] = 8'he5 ;
            rom[7747] = 8'h0b ;
            rom[7748] = 8'hfe ;
            rom[7749] = 8'hd5 ;
            rom[7750] = 8'h09 ;
            rom[7751] = 8'hfb ;
            rom[7752] = 8'hfb ;
            rom[7753] = 8'hee ;
            rom[7754] = 8'h18 ;
            rom[7755] = 8'h1b ;
            rom[7756] = 8'hff ;
            rom[7757] = 8'h17 ;
            rom[7758] = 8'hff ;
            rom[7759] = 8'h0a ;
            rom[7760] = 8'hb7 ;
            rom[7761] = 8'hf3 ;
            rom[7762] = 8'hd8 ;
            rom[7763] = 8'h0a ;
            rom[7764] = 8'h06 ;
            rom[7765] = 8'hfe ;
            rom[7766] = 8'h06 ;
            rom[7767] = 8'he8 ;
            rom[7768] = 8'h0e ;
            rom[7769] = 8'h11 ;
            rom[7770] = 8'h06 ;
            rom[7771] = 8'h14 ;
            rom[7772] = 8'h0d ;
            rom[7773] = 8'h0f ;
            rom[7774] = 8'h05 ;
            rom[7775] = 8'hfd ;
            rom[7776] = 8'hf5 ;
            rom[7777] = 8'hd4 ;
            rom[7778] = 8'h14 ;
            rom[7779] = 8'hf2 ;
            rom[7780] = 8'hd9 ;
            rom[7781] = 8'hb7 ;
            rom[7782] = 8'h14 ;
            rom[7783] = 8'h21 ;
            rom[7784] = 8'hdb ;
            rom[7785] = 8'he5 ;
            rom[7786] = 8'hf2 ;
            rom[7787] = 8'hf4 ;
            rom[7788] = 8'hcd ;
            rom[7789] = 8'h0c ;
            rom[7790] = 8'hf5 ;
            rom[7791] = 8'h1f ;
            rom[7792] = 8'h23 ;
            rom[7793] = 8'hef ;
            rom[7794] = 8'hfc ;
            rom[7795] = 8'h07 ;
            rom[7796] = 8'hed ;
            rom[7797] = 8'he8 ;
            rom[7798] = 8'hff ;
            rom[7799] = 8'hf7 ;
            rom[7800] = 8'hfe ;
            rom[7801] = 8'h17 ;
            rom[7802] = 8'h01 ;
            rom[7803] = 8'hf1 ;
            rom[7804] = 8'h07 ;
            rom[7805] = 8'h0a ;
            rom[7806] = 8'hdc ;
            rom[7807] = 8'h0d ;
            rom[7808] = 8'he9 ;
            rom[7809] = 8'hdd ;
            rom[7810] = 8'hf4 ;
            rom[7811] = 8'h0f ;
            rom[7812] = 8'hf8 ;
            rom[7813] = 8'hc4 ;
            rom[7814] = 8'h06 ;
            rom[7815] = 8'h27 ;
            rom[7816] = 8'hdd ;
            rom[7817] = 8'hfe ;
            rom[7818] = 8'hf9 ;
            rom[7819] = 8'hf4 ;
            rom[7820] = 8'he1 ;
            rom[7821] = 8'hea ;
            rom[7822] = 8'hfb ;
            rom[7823] = 8'hc6 ;
            rom[7824] = 8'hf3 ;
            rom[7825] = 8'he6 ;
            rom[7826] = 8'h16 ;
            rom[7827] = 8'hf7 ;
            rom[7828] = 8'h15 ;
            rom[7829] = 8'hde ;
            rom[7830] = 8'h0f ;
            rom[7831] = 8'hfd ;
            rom[7832] = 8'hdb ;
            rom[7833] = 8'h0d ;
            rom[7834] = 8'hf8 ;
            rom[7835] = 8'hf6 ;
            rom[7836] = 8'h1d ;
            rom[7837] = 8'h0b ;
            rom[7838] = 8'h0a ;
            rom[7839] = 8'h1c ;
            rom[7840] = 8'h13 ;
            rom[7841] = 8'h06 ;
            rom[7842] = 8'hf6 ;
            rom[7843] = 8'h2f ;
            rom[7844] = 8'h00 ;
            rom[7845] = 8'h06 ;
            rom[7846] = 8'hdd ;
            rom[7847] = 8'hfc ;
            rom[7848] = 8'hfa ;
            rom[7849] = 8'h0c ;
            rom[7850] = 8'hbf ;
            rom[7851] = 8'hf0 ;
            rom[7852] = 8'h05 ;
            rom[7853] = 8'he1 ;
            rom[7854] = 8'he6 ;
            rom[7855] = 8'h19 ;
            rom[7856] = 8'h0a ;
            rom[7857] = 8'hfa ;
            rom[7858] = 8'hf9 ;
            rom[7859] = 8'h15 ;
            rom[7860] = 8'he5 ;
            rom[7861] = 8'hef ;
            rom[7862] = 8'h01 ;
            rom[7863] = 8'hf1 ;
            rom[7864] = 8'hf3 ;
            rom[7865] = 8'h1b ;
            rom[7866] = 8'h15 ;
            rom[7867] = 8'heb ;
            rom[7868] = 8'hf4 ;
            rom[7869] = 8'hfd ;
            rom[7870] = 8'hf0 ;
            rom[7871] = 8'hf2 ;
            rom[7872] = 8'h09 ;
            rom[7873] = 8'h19 ;
            rom[7874] = 8'hff ;
            rom[7875] = 8'h9d ;
            rom[7876] = 8'hfc ;
            rom[7877] = 8'h08 ;
            rom[7878] = 8'hd5 ;
            rom[7879] = 8'hde ;
            rom[7880] = 8'h00 ;
            rom[7881] = 8'hf3 ;
            rom[7882] = 8'he2 ;
            rom[7883] = 8'hff ;
            rom[7884] = 8'hfa ;
            rom[7885] = 8'he3 ;
            rom[7886] = 8'hd8 ;
            rom[7887] = 8'h25 ;
            rom[7888] = 8'h0c ;
            rom[7889] = 8'hdd ;
            rom[7890] = 8'hf8 ;
            rom[7891] = 8'hd9 ;
            rom[7892] = 8'hfc ;
            rom[7893] = 8'he5 ;
            rom[7894] = 8'h09 ;
            rom[7895] = 8'hed ;
            rom[7896] = 8'h0b ;
            rom[7897] = 8'hf2 ;
            rom[7898] = 8'h1d ;
            rom[7899] = 8'h14 ;
            rom[7900] = 8'hf8 ;
            rom[7901] = 8'hfa ;
            rom[7902] = 8'h02 ;
            rom[7903] = 8'he9 ;
            rom[7904] = 8'hcd ;
            rom[7905] = 8'hff ;
            rom[7906] = 8'hf5 ;
            rom[7907] = 8'h05 ;
            rom[7908] = 8'hcf ;
            rom[7909] = 8'h0a ;
            rom[7910] = 8'hf1 ;
            rom[7911] = 8'hef ;
            rom[7912] = 8'he4 ;
            rom[7913] = 8'h06 ;
            rom[7914] = 8'h38 ;
            rom[7915] = 8'h08 ;
            rom[7916] = 8'hd9 ;
            rom[7917] = 8'h04 ;
            rom[7918] = 8'hec ;
            rom[7919] = 8'he2 ;
            rom[7920] = 8'h01 ;
            rom[7921] = 8'hff ;
            rom[7922] = 8'hd6 ;
            rom[7923] = 8'hee ;
            rom[7924] = 8'h15 ;
            rom[7925] = 8'hf7 ;
            rom[7926] = 8'hcb ;
            rom[7927] = 8'hf1 ;
            rom[7928] = 8'h08 ;
            rom[7929] = 8'hd4 ;
            rom[7930] = 8'hd9 ;
            rom[7931] = 8'h33 ;
            rom[7932] = 8'he6 ;
            rom[7933] = 8'he4 ;
            rom[7934] = 8'h10 ;
            rom[7935] = 8'he8 ;
            rom[7936] = 8'hcb ;
            rom[7937] = 8'h01 ;
            rom[7938] = 8'h09 ;
            rom[7939] = 8'h0e ;
            rom[7940] = 8'h09 ;
            rom[7941] = 8'h1b ;
            rom[7942] = 8'hea ;
            rom[7943] = 8'hfb ;
            rom[7944] = 8'hff ;
            rom[7945] = 8'h04 ;
            rom[7946] = 8'h05 ;
            rom[7947] = 8'hfa ;
            rom[7948] = 8'hd7 ;
            rom[7949] = 8'h18 ;
            rom[7950] = 8'h0e ;
            rom[7951] = 8'h19 ;
            rom[7952] = 8'h05 ;
            rom[7953] = 8'h1d ;
            rom[7954] = 8'he3 ;
            rom[7955] = 8'h0e ;
            rom[7956] = 8'h1d ;
            rom[7957] = 8'hf4 ;
            rom[7958] = 8'hef ;
            rom[7959] = 8'h11 ;
            rom[7960] = 8'hf1 ;
            rom[7961] = 8'h11 ;
            rom[7962] = 8'h00 ;
            rom[7963] = 8'he9 ;
            rom[7964] = 8'h07 ;
            rom[7965] = 8'hfe ;
            rom[7966] = 8'hed ;
            rom[7967] = 8'hf1 ;
            rom[7968] = 8'hea ;
            rom[7969] = 8'h28 ;
            rom[7970] = 8'h1b ;
            rom[7971] = 8'h1c ;
            rom[7972] = 8'hcf ;
            rom[7973] = 8'hfd ;
            rom[7974] = 8'hf3 ;
            rom[7975] = 8'hec ;
            rom[7976] = 8'h04 ;
            rom[7977] = 8'hf1 ;
            rom[7978] = 8'hf2 ;
            rom[7979] = 8'h14 ;
            rom[7980] = 8'heb ;
            rom[7981] = 8'hd5 ;
            rom[7982] = 8'h0e ;
            rom[7983] = 8'hcf ;
            rom[7984] = 8'hcf ;
            rom[7985] = 8'hce ;
            rom[7986] = 8'he8 ;
            rom[7987] = 8'hf3 ;
            rom[7988] = 8'h16 ;
            rom[7989] = 8'hee ;
            rom[7990] = 8'hf4 ;
            rom[7991] = 8'hcc ;
            rom[7992] = 8'hfe ;
            rom[7993] = 8'he7 ;
            rom[7994] = 8'hfa ;
            rom[7995] = 8'hd1 ;
            rom[7996] = 8'he3 ;
            rom[7997] = 8'hd1 ;
            rom[7998] = 8'h10 ;
            rom[7999] = 8'h14 ;
            rom[8000] = 8'hf8 ;
            rom[8001] = 8'hee ;
            rom[8002] = 8'hd3 ;
            rom[8003] = 8'h08 ;
            rom[8004] = 8'hf8 ;
            rom[8005] = 8'hd7 ;
            rom[8006] = 8'hd7 ;
            rom[8007] = 8'h2a ;
            rom[8008] = 8'hd4 ;
            rom[8009] = 8'hf4 ;
            rom[8010] = 8'h21 ;
            rom[8011] = 8'h01 ;
            rom[8012] = 8'h0d ;
            rom[8013] = 8'h13 ;
            rom[8014] = 8'h26 ;
            rom[8015] = 8'h15 ;
            rom[8016] = 8'hf8 ;
            rom[8017] = 8'hf8 ;
            rom[8018] = 8'h03 ;
            rom[8019] = 8'h0e ;
            rom[8020] = 8'h16 ;
            rom[8021] = 8'hf2 ;
            rom[8022] = 8'hfe ;
            rom[8023] = 8'h0a ;
            rom[8024] = 8'h1d ;
            rom[8025] = 8'hf9 ;
            rom[8026] = 8'hf6 ;
            rom[8027] = 8'hf2 ;
            rom[8028] = 8'hf2 ;
            rom[8029] = 8'h0d ;
            rom[8030] = 8'hfa ;
            rom[8031] = 8'h17 ;
            rom[8032] = 8'hf5 ;
            rom[8033] = 8'h07 ;
            rom[8034] = 8'h10 ;
            rom[8035] = 8'hc1 ;
            rom[8036] = 8'he0 ;
            rom[8037] = 8'hc4 ;
            rom[8038] = 8'hf4 ;
            rom[8039] = 8'h2f ;
            rom[8040] = 8'hfb ;
            rom[8041] = 8'h11 ;
            rom[8042] = 8'hc0 ;
            rom[8043] = 8'hf9 ;
            rom[8044] = 8'h0c ;
            rom[8045] = 8'he2 ;
            rom[8046] = 8'hf4 ;
            rom[8047] = 8'h1c ;
            rom[8048] = 8'h15 ;
            rom[8049] = 8'h1e ;
            rom[8050] = 8'h06 ;
            rom[8051] = 8'h19 ;
            rom[8052] = 8'h12 ;
            rom[8053] = 8'hfb ;
            rom[8054] = 8'h1f ;
            rom[8055] = 8'h09 ;
            rom[8056] = 8'h09 ;
            rom[8057] = 8'h1a ;
            rom[8058] = 8'h0f ;
            rom[8059] = 8'hd4 ;
            rom[8060] = 8'h22 ;
            rom[8061] = 8'h04 ;
            rom[8062] = 8'hd2 ;
            rom[8063] = 8'h00 ;
            rom[8064] = 8'h0c ;
            rom[8065] = 8'h19 ;
            rom[8066] = 8'h08 ;
            rom[8067] = 8'hd6 ;
            rom[8068] = 8'hf0 ;
            rom[8069] = 8'he8 ;
            rom[8070] = 8'h35 ;
            rom[8071] = 8'h07 ;
            rom[8072] = 8'hf9 ;
            rom[8073] = 8'h01 ;
            rom[8074] = 8'hde ;
            rom[8075] = 8'hf9 ;
            rom[8076] = 8'h12 ;
            rom[8077] = 8'hed ;
            rom[8078] = 8'h28 ;
            rom[8079] = 8'h04 ;
            rom[8080] = 8'h0b ;
            rom[8081] = 8'hf1 ;
            rom[8082] = 8'h1a ;
            rom[8083] = 8'h1d ;
            rom[8084] = 8'hee ;
            rom[8085] = 8'hcd ;
            rom[8086] = 8'hc8 ;
            rom[8087] = 8'he4 ;
            rom[8088] = 8'hd7 ;
            rom[8089] = 8'hf8 ;
            rom[8090] = 8'hc7 ;
            rom[8091] = 8'hbd ;
            rom[8092] = 8'h09 ;
            rom[8093] = 8'hfe ;
            rom[8094] = 8'hd4 ;
            rom[8095] = 8'hec ;
            rom[8096] = 8'hc4 ;
            rom[8097] = 8'hef ;
            rom[8098] = 8'h21 ;
            rom[8099] = 8'h12 ;
            rom[8100] = 8'h03 ;
            rom[8101] = 8'hda ;
            rom[8102] = 8'h08 ;
            rom[8103] = 8'hcd ;
            rom[8104] = 8'h05 ;
            rom[8105] = 8'h07 ;
            rom[8106] = 8'hf7 ;
            rom[8107] = 8'hf3 ;
            rom[8108] = 8'h0c ;
            rom[8109] = 8'hf4 ;
            rom[8110] = 8'h0e ;
            rom[8111] = 8'hca ;
            rom[8112] = 8'hf6 ;
            rom[8113] = 8'hc7 ;
            rom[8114] = 8'hdf ;
            rom[8115] = 8'h07 ;
            rom[8116] = 8'hdc ;
            rom[8117] = 8'h17 ;
            rom[8118] = 8'hfd ;
            rom[8119] = 8'hf7 ;
            rom[8120] = 8'he5 ;
            rom[8121] = 8'hf9 ;
            rom[8122] = 8'hdf ;
            rom[8123] = 8'hef ;
            rom[8124] = 8'hcd ;
            rom[8125] = 8'hc0 ;
            rom[8126] = 8'hfc ;
            rom[8127] = 8'h10 ;
            rom[8128] = 8'h17 ;
            rom[8129] = 8'h0f ;
            rom[8130] = 8'he2 ;
            rom[8131] = 8'hd3 ;
            rom[8132] = 8'hdc ;
            rom[8133] = 8'h0c ;
            rom[8134] = 8'h00 ;
            rom[8135] = 8'hf7 ;
            rom[8136] = 8'hf8 ;
            rom[8137] = 8'h07 ;
            rom[8138] = 8'h0e ;
            rom[8139] = 8'h20 ;
            rom[8140] = 8'h01 ;
            rom[8141] = 8'hdc ;
            rom[8142] = 8'h0f ;
            rom[8143] = 8'hc7 ;
            rom[8144] = 8'h0a ;
            rom[8145] = 8'hbe ;
            rom[8146] = 8'hde ;
            rom[8147] = 8'hf1 ;
            rom[8148] = 8'h2a ;
            rom[8149] = 8'h0c ;
            rom[8150] = 8'hed ;
            rom[8151] = 8'h02 ;
            rom[8152] = 8'hea ;
            rom[8153] = 8'hdc ;
            rom[8154] = 8'h08 ;
            rom[8155] = 8'hf3 ;
            rom[8156] = 8'hc7 ;
            rom[8157] = 8'hc8 ;
            rom[8158] = 8'hd8 ;
            rom[8159] = 8'hea ;
            rom[8160] = 8'hef ;
            rom[8161] = 8'hf4 ;
            rom[8162] = 8'h18 ;
            rom[8163] = 8'hfb ;
            rom[8164] = 8'hf6 ;
            rom[8165] = 8'hfe ;
            rom[8166] = 8'hf5 ;
            rom[8167] = 8'hfa ;
            rom[8168] = 8'h02 ;
            rom[8169] = 8'hf6 ;
            rom[8170] = 8'hf7 ;
            rom[8171] = 8'he2 ;
            rom[8172] = 8'h0c ;
            rom[8173] = 8'hef ;
            rom[8174] = 8'h11 ;
            rom[8175] = 8'hfc ;
            rom[8176] = 8'hed ;
            rom[8177] = 8'h02 ;
            rom[8178] = 8'h13 ;
            rom[8179] = 8'hd8 ;
            rom[8180] = 8'h10 ;
            rom[8181] = 8'h28 ;
            rom[8182] = 8'h06 ;
            rom[8183] = 8'h18 ;
            rom[8184] = 8'hda ;
            rom[8185] = 8'hd2 ;
            rom[8186] = 8'hf5 ;
            rom[8187] = 8'hc5 ;
            rom[8188] = 8'hfa ;
            rom[8189] = 8'hc4 ;
            rom[8190] = 8'hfe ;
            rom[8191] = 8'h0b ;
            rom[8192] = 8'hff ;
            rom[8193] = 8'hee ;
            rom[8194] = 8'h00 ;
            rom[8195] = 8'hf3 ;
            rom[8196] = 8'hee ;
            rom[8197] = 8'hfe ;
            rom[8198] = 8'h11 ;
            rom[8199] = 8'hc2 ;
            rom[8200] = 8'h02 ;
            rom[8201] = 8'h03 ;
            rom[8202] = 8'h0b ;
            rom[8203] = 8'h05 ;
            rom[8204] = 8'h1d ;
            rom[8205] = 8'hda ;
            rom[8206] = 8'h14 ;
            rom[8207] = 8'h07 ;
            rom[8208] = 8'hea ;
            rom[8209] = 8'hd3 ;
            rom[8210] = 8'hee ;
            rom[8211] = 8'he3 ;
            rom[8212] = 8'h13 ;
            rom[8213] = 8'h20 ;
            rom[8214] = 8'h0a ;
            rom[8215] = 8'he7 ;
            rom[8216] = 8'h0a ;
            rom[8217] = 8'he6 ;
            rom[8218] = 8'heb ;
            rom[8219] = 8'h19 ;
            rom[8220] = 8'hf7 ;
            rom[8221] = 8'hff ;
            rom[8222] = 8'h05 ;
            rom[8223] = 8'h11 ;
            rom[8224] = 8'hf4 ;
            rom[8225] = 8'he8 ;
            rom[8226] = 8'hec ;
            rom[8227] = 8'hf4 ;
            rom[8228] = 8'h2f ;
            rom[8229] = 8'h16 ;
            rom[8230] = 8'h10 ;
            rom[8231] = 8'h05 ;
            rom[8232] = 8'hfc ;
            rom[8233] = 8'he3 ;
            rom[8234] = 8'h0d ;
            rom[8235] = 8'hf3 ;
            rom[8236] = 8'h0b ;
            rom[8237] = 8'h06 ;
            rom[8238] = 8'hf2 ;
            rom[8239] = 8'hcb ;
            rom[8240] = 8'hf7 ;
            rom[8241] = 8'h08 ;
            rom[8242] = 8'hd0 ;
            rom[8243] = 8'h0e ;
            rom[8244] = 8'hf6 ;
            rom[8245] = 8'h19 ;
            rom[8246] = 8'hc0 ;
            rom[8247] = 8'hcc ;
            rom[8248] = 8'h12 ;
            rom[8249] = 8'he7 ;
            rom[8250] = 8'hf8 ;
            rom[8251] = 8'h23 ;
            rom[8252] = 8'h08 ;
            rom[8253] = 8'hfc ;
            rom[8254] = 8'h0c ;
            rom[8255] = 8'hce ;
            rom[8256] = 8'he9 ;
            rom[8257] = 8'h0e ;
            rom[8258] = 8'h0c ;
            rom[8259] = 8'h0f ;
            rom[8260] = 8'hfe ;
            rom[8261] = 8'h04 ;
            rom[8262] = 8'h02 ;
            rom[8263] = 8'h12 ;
            rom[8264] = 8'h00 ;
            rom[8265] = 8'h0d ;
            rom[8266] = 8'hf2 ;
            rom[8267] = 8'h0b ;
            rom[8268] = 8'hf9 ;
            rom[8269] = 8'hd9 ;
            rom[8270] = 8'he1 ;
            rom[8271] = 8'he3 ;
            rom[8272] = 8'h1a ;
            rom[8273] = 8'h07 ;
            rom[8274] = 8'h11 ;
            rom[8275] = 8'h0d ;
            rom[8276] = 8'he9 ;
            rom[8277] = 8'hdd ;
            rom[8278] = 8'h03 ;
            rom[8279] = 8'hd0 ;
            rom[8280] = 8'h11 ;
            rom[8281] = 8'hf8 ;
            rom[8282] = 8'h0f ;
            rom[8283] = 8'h06 ;
            rom[8284] = 8'hf8 ;
            rom[8285] = 8'h0f ;
            rom[8286] = 8'he8 ;
            rom[8287] = 8'h07 ;
            rom[8288] = 8'hf3 ;
            rom[8289] = 8'h1f ;
            rom[8290] = 8'hd9 ;
            rom[8291] = 8'hce ;
            rom[8292] = 8'h0a ;
            rom[8293] = 8'hfc ;
            rom[8294] = 8'h26 ;
            rom[8295] = 8'h0a ;
            rom[8296] = 8'hf3 ;
            rom[8297] = 8'h18 ;
            rom[8298] = 8'hf5 ;
            rom[8299] = 8'h08 ;
            rom[8300] = 8'hf1 ;
            rom[8301] = 8'h02 ;
            rom[8302] = 8'h03 ;
            rom[8303] = 8'h1d ;
            rom[8304] = 8'h12 ;
            rom[8305] = 8'hcf ;
            rom[8306] = 8'h04 ;
            rom[8307] = 8'h07 ;
            rom[8308] = 8'h0f ;
            rom[8309] = 8'h11 ;
            rom[8310] = 8'hf0 ;
            rom[8311] = 8'hd7 ;
            rom[8312] = 8'h03 ;
            rom[8313] = 8'h0e ;
            rom[8314] = 8'h1b ;
            rom[8315] = 8'hf3 ;
            rom[8316] = 8'hf7 ;
            rom[8317] = 8'hd9 ;
            rom[8318] = 8'he5 ;
            rom[8319] = 8'hf1 ;
            rom[8320] = 8'h0f ;
            rom[8321] = 8'h03 ;
            rom[8322] = 8'h15 ;
            rom[8323] = 8'h00 ;
            rom[8324] = 8'hfb ;
            rom[8325] = 8'he2 ;
            rom[8326] = 8'hea ;
            rom[8327] = 8'he7 ;
            rom[8328] = 8'hfc ;
            rom[8329] = 8'hf5 ;
            rom[8330] = 8'h0f ;
            rom[8331] = 8'h02 ;
            rom[8332] = 8'h02 ;
            rom[8333] = 8'hf8 ;
            rom[8334] = 8'hec ;
            rom[8335] = 8'hd3 ;
            rom[8336] = 8'hea ;
            rom[8337] = 8'hfe ;
            rom[8338] = 8'h21 ;
            rom[8339] = 8'hef ;
            rom[8340] = 8'he8 ;
            rom[8341] = 8'hc3 ;
            rom[8342] = 8'h1b ;
            rom[8343] = 8'hf2 ;
            rom[8344] = 8'hda ;
            rom[8345] = 8'hef ;
            rom[8346] = 8'hef ;
            rom[8347] = 8'hd0 ;
            rom[8348] = 8'h07 ;
            rom[8349] = 8'hd5 ;
            rom[8350] = 8'hf6 ;
            rom[8351] = 8'heb ;
            rom[8352] = 8'hd3 ;
            rom[8353] = 8'h19 ;
            rom[8354] = 8'hd4 ;
            rom[8355] = 8'h1d ;
            rom[8356] = 8'hde ;
            rom[8357] = 8'hf0 ;
            rom[8358] = 8'hee ;
            rom[8359] = 8'hec ;
            rom[8360] = 8'hfb ;
            rom[8361] = 8'heb ;
            rom[8362] = 8'h00 ;
            rom[8363] = 8'he4 ;
            rom[8364] = 8'hb7 ;
            rom[8365] = 8'he0 ;
            rom[8366] = 8'hf1 ;
            rom[8367] = 8'h09 ;
            rom[8368] = 8'he3 ;
            rom[8369] = 8'hf8 ;
            rom[8370] = 8'hea ;
            rom[8371] = 8'h0e ;
            rom[8372] = 8'h03 ;
            rom[8373] = 8'hfb ;
            rom[8374] = 8'hd6 ;
            rom[8375] = 8'hfc ;
            rom[8376] = 8'hf9 ;
            rom[8377] = 8'hf0 ;
            rom[8378] = 8'he0 ;
            rom[8379] = 8'h0d ;
            rom[8380] = 8'hd3 ;
            rom[8381] = 8'hfa ;
            rom[8382] = 8'hcf ;
            rom[8383] = 8'hdd ;
            rom[8384] = 8'h03 ;
            rom[8385] = 8'he4 ;
            rom[8386] = 8'hf4 ;
            rom[8387] = 8'hed ;
            rom[8388] = 8'hf9 ;
            rom[8389] = 8'hd7 ;
            rom[8390] = 8'hed ;
            rom[8391] = 8'he5 ;
            rom[8392] = 8'h03 ;
            rom[8393] = 8'h11 ;
            rom[8394] = 8'h12 ;
            rom[8395] = 8'h00 ;
            rom[8396] = 8'hec ;
            rom[8397] = 8'h0d ;
            rom[8398] = 8'h11 ;
            rom[8399] = 8'h08 ;
            rom[8400] = 8'hf3 ;
            rom[8401] = 8'hfc ;
            rom[8402] = 8'hd9 ;
            rom[8403] = 8'h07 ;
            rom[8404] = 8'hf8 ;
            rom[8405] = 8'hc3 ;
            rom[8406] = 8'h05 ;
            rom[8407] = 8'hef ;
            rom[8408] = 8'h03 ;
            rom[8409] = 8'h01 ;
            rom[8410] = 8'h04 ;
            rom[8411] = 8'he6 ;
            rom[8412] = 8'hcd ;
            rom[8413] = 8'hd9 ;
            rom[8414] = 8'hff ;
            rom[8415] = 8'hfc ;
            rom[8416] = 8'hdd ;
            rom[8417] = 8'hf3 ;
            rom[8418] = 8'hfa ;
            rom[8419] = 8'hdf ;
            rom[8420] = 8'h04 ;
            rom[8421] = 8'hfa ;
            rom[8422] = 8'hde ;
            rom[8423] = 8'hf7 ;
            rom[8424] = 8'hd0 ;
            rom[8425] = 8'he6 ;
            rom[8426] = 8'hd4 ;
            rom[8427] = 8'hec ;
            rom[8428] = 8'hee ;
            rom[8429] = 8'hfb ;
            rom[8430] = 8'h14 ;
            rom[8431] = 8'h15 ;
            rom[8432] = 8'hec ;
            rom[8433] = 8'hf2 ;
            rom[8434] = 8'h0a ;
            rom[8435] = 8'hf5 ;
            rom[8436] = 8'hb1 ;
            rom[8437] = 8'h20 ;
            rom[8438] = 8'h0e ;
            rom[8439] = 8'hef ;
            rom[8440] = 8'hf7 ;
            rom[8441] = 8'h21 ;
            rom[8442] = 8'h10 ;
            rom[8443] = 8'hfb ;
            rom[8444] = 8'h09 ;
            rom[8445] = 8'haf ;
            rom[8446] = 8'hc6 ;
            rom[8447] = 8'hd1 ;
            rom[8448] = 8'h04 ;
            rom[8449] = 8'he1 ;
            rom[8450] = 8'he5 ;
            rom[8451] = 8'hfd ;
            rom[8452] = 8'hf5 ;
            rom[8453] = 8'hed ;
            rom[8454] = 8'h02 ;
            rom[8455] = 8'hc7 ;
            rom[8456] = 8'h01 ;
            rom[8457] = 8'h0b ;
            rom[8458] = 8'hd5 ;
            rom[8459] = 8'h02 ;
            rom[8460] = 8'hdb ;
            rom[8461] = 8'hfc ;
            rom[8462] = 8'h06 ;
            rom[8463] = 8'h01 ;
            rom[8464] = 8'h06 ;
            rom[8465] = 8'h15 ;
            rom[8466] = 8'hd0 ;
            rom[8467] = 8'hfd ;
            rom[8468] = 8'h20 ;
            rom[8469] = 8'h0d ;
            rom[8470] = 8'hcc ;
            rom[8471] = 8'hf1 ;
            rom[8472] = 8'h04 ;
            rom[8473] = 8'h24 ;
            rom[8474] = 8'h0c ;
            rom[8475] = 8'hfa ;
            rom[8476] = 8'h1a ;
            rom[8477] = 8'h2b ;
            rom[8478] = 8'hf6 ;
            rom[8479] = 8'hf7 ;
            rom[8480] = 8'h1a ;
            rom[8481] = 8'hf3 ;
            rom[8482] = 8'h1f ;
            rom[8483] = 8'he6 ;
            rom[8484] = 8'hd1 ;
            rom[8485] = 8'hdd ;
            rom[8486] = 8'heb ;
            rom[8487] = 8'hf8 ;
            rom[8488] = 8'he3 ;
            rom[8489] = 8'h07 ;
            rom[8490] = 8'hda ;
            rom[8491] = 8'hc9 ;
            rom[8492] = 8'h1b ;
            rom[8493] = 8'h24 ;
            rom[8494] = 8'h07 ;
            rom[8495] = 8'hef ;
            rom[8496] = 8'hd7 ;
            rom[8497] = 8'h11 ;
            rom[8498] = 8'he9 ;
            rom[8499] = 8'hc9 ;
            rom[8500] = 8'h10 ;
            rom[8501] = 8'hff ;
            rom[8502] = 8'ha6 ;
            rom[8503] = 8'hf2 ;
            rom[8504] = 8'h10 ;
            rom[8505] = 8'h0a ;
            rom[8506] = 8'hfe ;
            rom[8507] = 8'hc7 ;
            rom[8508] = 8'heb ;
            rom[8509] = 8'hae ;
            rom[8510] = 8'hf3 ;
            rom[8511] = 8'hfb ;
            rom[8512] = 8'h02 ;
            rom[8513] = 8'h09 ;
            rom[8514] = 8'h03 ;
            rom[8515] = 8'h16 ;
            rom[8516] = 8'h05 ;
            rom[8517] = 8'heb ;
            rom[8518] = 8'hf9 ;
            rom[8519] = 8'h0d ;
            rom[8520] = 8'he6 ;
            rom[8521] = 8'hf1 ;
            rom[8522] = 8'h14 ;
            rom[8523] = 8'h1f ;
            rom[8524] = 8'h17 ;
            rom[8525] = 8'hff ;
            rom[8526] = 8'hfc ;
            rom[8527] = 8'h2f ;
            rom[8528] = 8'hf4 ;
            rom[8529] = 8'hda ;
            rom[8530] = 8'hf8 ;
            rom[8531] = 8'h0f ;
            rom[8532] = 8'hf4 ;
            rom[8533] = 8'h23 ;
            rom[8534] = 8'hcd ;
            rom[8535] = 8'hfa ;
            rom[8536] = 8'h0c ;
            rom[8537] = 8'hf9 ;
            rom[8538] = 8'hfa ;
            rom[8539] = 8'h17 ;
            rom[8540] = 8'h1c ;
            rom[8541] = 8'h1f ;
            rom[8542] = 8'h18 ;
            rom[8543] = 8'hf4 ;
            rom[8544] = 8'h11 ;
            rom[8545] = 8'he4 ;
            rom[8546] = 8'h15 ;
            rom[8547] = 8'hcf ;
            rom[8548] = 8'hce ;
            rom[8549] = 8'h0b ;
            rom[8550] = 8'he7 ;
            rom[8551] = 8'h12 ;
            rom[8552] = 8'hef ;
            rom[8553] = 8'hd4 ;
            rom[8554] = 8'h1a ;
            rom[8555] = 8'hf6 ;
            rom[8556] = 8'h13 ;
            rom[8557] = 8'h07 ;
            rom[8558] = 8'hf7 ;
            rom[8559] = 8'h13 ;
            rom[8560] = 8'h02 ;
            rom[8561] = 8'h01 ;
            rom[8562] = 8'h06 ;
            rom[8563] = 8'hf8 ;
            rom[8564] = 8'h0e ;
            rom[8565] = 8'hf5 ;
            rom[8566] = 8'h08 ;
            rom[8567] = 8'hf5 ;
            rom[8568] = 8'hf7 ;
            rom[8569] = 8'hdb ;
            rom[8570] = 8'hf1 ;
            rom[8571] = 8'hef ;
            rom[8572] = 8'h02 ;
            rom[8573] = 8'heb ;
            rom[8574] = 8'he5 ;
            rom[8575] = 8'hf2 ;
            rom[8576] = 8'h9e ;
            rom[8577] = 8'h0d ;
            rom[8578] = 8'h15 ;
            rom[8579] = 8'h03 ;
            rom[8580] = 8'h0d ;
            rom[8581] = 8'he9 ;
            rom[8582] = 8'h1c ;
            rom[8583] = 8'h01 ;
            rom[8584] = 8'hda ;
            rom[8585] = 8'hf0 ;
            rom[8586] = 8'hf4 ;
            rom[8587] = 8'hf4 ;
            rom[8588] = 8'hf1 ;
            rom[8589] = 8'h13 ;
            rom[8590] = 8'h09 ;
            rom[8591] = 8'h08 ;
            rom[8592] = 8'h02 ;
            rom[8593] = 8'hcf ;
            rom[8594] = 8'he0 ;
            rom[8595] = 8'hda ;
            rom[8596] = 8'h17 ;
            rom[8597] = 8'h02 ;
            rom[8598] = 8'hea ;
            rom[8599] = 8'hf7 ;
            rom[8600] = 8'hfc ;
            rom[8601] = 8'hfb ;
            rom[8602] = 8'h0e ;
            rom[8603] = 8'hec ;
            rom[8604] = 8'h0a ;
            rom[8605] = 8'h07 ;
            rom[8606] = 8'he8 ;
            rom[8607] = 8'hd7 ;
            rom[8608] = 8'h0d ;
            rom[8609] = 8'hd5 ;
            rom[8610] = 8'h09 ;
            rom[8611] = 8'h0b ;
            rom[8612] = 8'h1e ;
            rom[8613] = 8'h02 ;
            rom[8614] = 8'h0c ;
            rom[8615] = 8'h12 ;
            rom[8616] = 8'hff ;
            rom[8617] = 8'hdd ;
            rom[8618] = 8'hfd ;
            rom[8619] = 8'hef ;
            rom[8620] = 8'h06 ;
            rom[8621] = 8'hf5 ;
            rom[8622] = 8'h0c ;
            rom[8623] = 8'hde ;
            rom[8624] = 8'h36 ;
            rom[8625] = 8'h09 ;
            rom[8626] = 8'hfd ;
            rom[8627] = 8'hde ;
            rom[8628] = 8'hed ;
            rom[8629] = 8'h19 ;
            rom[8630] = 8'hfa ;
            rom[8631] = 8'he3 ;
            rom[8632] = 8'hde ;
            rom[8633] = 8'hf7 ;
            rom[8634] = 8'hfa ;
            rom[8635] = 8'hfe ;
            rom[8636] = 8'he9 ;
            rom[8637] = 8'hf8 ;
            rom[8638] = 8'h08 ;
            rom[8639] = 8'he2 ;
            rom[8640] = 8'he9 ;
            rom[8641] = 8'hff ;
            rom[8642] = 8'he7 ;
            rom[8643] = 8'h07 ;
            rom[8644] = 8'hdb ;
            rom[8645] = 8'hd7 ;
            rom[8646] = 8'hfc ;
            rom[8647] = 8'h16 ;
            rom[8648] = 8'hbf ;
            rom[8649] = 8'hee ;
            rom[8650] = 8'hf8 ;
            rom[8651] = 8'h2b ;
            rom[8652] = 8'h0e ;
            rom[8653] = 8'hdf ;
            rom[8654] = 8'he0 ;
            rom[8655] = 8'h17 ;
            rom[8656] = 8'hf4 ;
            rom[8657] = 8'hf9 ;
            rom[8658] = 8'he8 ;
            rom[8659] = 8'h07 ;
            rom[8660] = 8'he0 ;
            rom[8661] = 8'h16 ;
            rom[8662] = 8'hf6 ;
            rom[8663] = 8'he6 ;
            rom[8664] = 8'h2e ;
            rom[8665] = 8'hfb ;
            rom[8666] = 8'h1d ;
            rom[8667] = 8'h0a ;
            rom[8668] = 8'hf1 ;
            rom[8669] = 8'h13 ;
            rom[8670] = 8'hd1 ;
            rom[8671] = 8'h09 ;
            rom[8672] = 8'he7 ;
            rom[8673] = 8'h15 ;
            rom[8674] = 8'hfe ;
            rom[8675] = 8'hfe ;
            rom[8676] = 8'h22 ;
            rom[8677] = 8'hff ;
            rom[8678] = 8'h2c ;
            rom[8679] = 8'h1f ;
            rom[8680] = 8'h03 ;
            rom[8681] = 8'hea ;
            rom[8682] = 8'h1d ;
            rom[8683] = 8'hf6 ;
            rom[8684] = 8'hfe ;
            rom[8685] = 8'he5 ;
            rom[8686] = 8'hd0 ;
            rom[8687] = 8'h0d ;
            rom[8688] = 8'h13 ;
            rom[8689] = 8'hee ;
            rom[8690] = 8'h1e ;
            rom[8691] = 8'h01 ;
            rom[8692] = 8'h0d ;
            rom[8693] = 8'h20 ;
            rom[8694] = 8'hec ;
            rom[8695] = 8'h0b ;
            rom[8696] = 8'h08 ;
            rom[8697] = 8'hf8 ;
            rom[8698] = 8'h17 ;
            rom[8699] = 8'h06 ;
            rom[8700] = 8'h1b ;
            rom[8701] = 8'h07 ;
            rom[8702] = 8'hfe ;
            rom[8703] = 8'h0a ;
            rom[8704] = 8'hfa ;
            rom[8705] = 8'h09 ;
            rom[8706] = 8'h1b ;
            rom[8707] = 8'h13 ;
            rom[8708] = 8'h07 ;
            rom[8709] = 8'h02 ;
            rom[8710] = 8'h14 ;
            rom[8711] = 8'hf1 ;
            rom[8712] = 8'h0b ;
            rom[8713] = 8'hf7 ;
            rom[8714] = 8'hed ;
            rom[8715] = 8'he2 ;
            rom[8716] = 8'h19 ;
            rom[8717] = 8'h0e ;
            rom[8718] = 8'hff ;
            rom[8719] = 8'hd7 ;
            rom[8720] = 8'hcc ;
            rom[8721] = 8'h10 ;
            rom[8722] = 8'h12 ;
            rom[8723] = 8'hf2 ;
            rom[8724] = 8'hf3 ;
            rom[8725] = 8'h14 ;
            rom[8726] = 8'h0d ;
            rom[8727] = 8'h12 ;
            rom[8728] = 8'hf0 ;
            rom[8729] = 8'hfc ;
            rom[8730] = 8'he2 ;
            rom[8731] = 8'h02 ;
            rom[8732] = 8'hfa ;
            rom[8733] = 8'he0 ;
            rom[8734] = 8'h0c ;
            rom[8735] = 8'h0c ;
            rom[8736] = 8'h0f ;
            rom[8737] = 8'h0a ;
            rom[8738] = 8'he9 ;
            rom[8739] = 8'hd4 ;
            rom[8740] = 8'hed ;
            rom[8741] = 8'hd2 ;
            rom[8742] = 8'h08 ;
            rom[8743] = 8'hf2 ;
            rom[8744] = 8'hea ;
            rom[8745] = 8'hf0 ;
            rom[8746] = 8'h04 ;
            rom[8747] = 8'h2e ;
            rom[8748] = 8'h12 ;
            rom[8749] = 8'hf7 ;
            rom[8750] = 8'he2 ;
            rom[8751] = 8'hff ;
            rom[8752] = 8'hd9 ;
            rom[8753] = 8'h10 ;
            rom[8754] = 8'h1d ;
            rom[8755] = 8'he7 ;
            rom[8756] = 8'h00 ;
            rom[8757] = 8'h0b ;
            rom[8758] = 8'h08 ;
            rom[8759] = 8'hfe ;
            rom[8760] = 8'h09 ;
            rom[8761] = 8'heb ;
            rom[8762] = 8'h1a ;
            rom[8763] = 8'hef ;
            rom[8764] = 8'hf7 ;
            rom[8765] = 8'h00 ;
            rom[8766] = 8'h11 ;
            rom[8767] = 8'hec ;
            rom[8768] = 8'h19 ;
            rom[8769] = 8'hee ;
            rom[8770] = 8'hea ;
            rom[8771] = 8'h16 ;
            rom[8772] = 8'h1b ;
            rom[8773] = 8'hf5 ;
            rom[8774] = 8'hdc ;
            rom[8775] = 8'hf6 ;
            rom[8776] = 8'hef ;
            rom[8777] = 8'hfb ;
            rom[8778] = 8'he3 ;
            rom[8779] = 8'he5 ;
            rom[8780] = 8'he8 ;
            rom[8781] = 8'h1a ;
            rom[8782] = 8'hc0 ;
            rom[8783] = 8'h08 ;
            rom[8784] = 8'hea ;
            rom[8785] = 8'h17 ;
            rom[8786] = 8'hee ;
            rom[8787] = 8'h09 ;
            rom[8788] = 8'hf6 ;
            rom[8789] = 8'hef ;
            rom[8790] = 8'hff ;
            rom[8791] = 8'hef ;
            rom[8792] = 8'he7 ;
            rom[8793] = 8'he5 ;
            rom[8794] = 8'hf3 ;
            rom[8795] = 8'hd1 ;
            rom[8796] = 8'hf2 ;
            rom[8797] = 8'hfb ;
            rom[8798] = 8'h11 ;
            rom[8799] = 8'he6 ;
            rom[8800] = 8'h16 ;
            rom[8801] = 8'h11 ;
            rom[8802] = 8'hc1 ;
            rom[8803] = 8'hfc ;
            rom[8804] = 8'hf7 ;
            rom[8805] = 8'he6 ;
            rom[8806] = 8'h05 ;
            rom[8807] = 8'hd7 ;
            rom[8808] = 8'hf7 ;
            rom[8809] = 8'hff ;
            rom[8810] = 8'hf9 ;
            rom[8811] = 8'h2b ;
            rom[8812] = 8'he5 ;
            rom[8813] = 8'h03 ;
            rom[8814] = 8'h03 ;
            rom[8815] = 8'h17 ;
            rom[8816] = 8'hef ;
            rom[8817] = 8'h0d ;
            rom[8818] = 8'hfb ;
            rom[8819] = 8'h15 ;
            rom[8820] = 8'hf1 ;
            rom[8821] = 8'hdb ;
            rom[8822] = 8'hf1 ;
            rom[8823] = 8'hff ;
            rom[8824] = 8'he5 ;
            rom[8825] = 8'he2 ;
            rom[8826] = 8'hc2 ;
            rom[8827] = 8'hf5 ;
            rom[8828] = 8'he8 ;
            rom[8829] = 8'h2c ;
            rom[8830] = 8'hf3 ;
            rom[8831] = 8'he1 ;
            rom[8832] = 8'hf6 ;
            rom[8833] = 8'he5 ;
            rom[8834] = 8'he3 ;
            rom[8835] = 8'h08 ;
            rom[8836] = 8'h22 ;
            rom[8837] = 8'he1 ;
            rom[8838] = 8'hd1 ;
            rom[8839] = 8'hfc ;
            rom[8840] = 8'hf5 ;
            rom[8841] = 8'h0f ;
            rom[8842] = 8'hf9 ;
            rom[8843] = 8'hf3 ;
            rom[8844] = 8'hdb ;
            rom[8845] = 8'hfc ;
            rom[8846] = 8'hfb ;
            rom[8847] = 8'he1 ;
            rom[8848] = 8'h1c ;
            rom[8849] = 8'h04 ;
            rom[8850] = 8'hfb ;
            rom[8851] = 8'hf5 ;
            rom[8852] = 8'h0b ;
            rom[8853] = 8'he8 ;
            rom[8854] = 8'hf4 ;
            rom[8855] = 8'h06 ;
            rom[8856] = 8'h08 ;
            rom[8857] = 8'hfd ;
            rom[8858] = 8'h1b ;
            rom[8859] = 8'h03 ;
            rom[8860] = 8'h00 ;
            rom[8861] = 8'h1a ;
            rom[8862] = 8'hfa ;
            rom[8863] = 8'h23 ;
            rom[8864] = 8'h11 ;
            rom[8865] = 8'h00 ;
            rom[8866] = 8'hca ;
            rom[8867] = 8'hf5 ;
            rom[8868] = 8'heb ;
            rom[8869] = 8'h06 ;
            rom[8870] = 8'hf8 ;
            rom[8871] = 8'h18 ;
            rom[8872] = 8'h27 ;
            rom[8873] = 8'hfb ;
            rom[8874] = 8'heb ;
            rom[8875] = 8'h02 ;
            rom[8876] = 8'he4 ;
            rom[8877] = 8'h02 ;
            rom[8878] = 8'hf0 ;
            rom[8879] = 8'h08 ;
            rom[8880] = 8'hf2 ;
            rom[8881] = 8'h1d ;
            rom[8882] = 8'h09 ;
            rom[8883] = 8'hee ;
            rom[8884] = 8'h21 ;
            rom[8885] = 8'hee ;
            rom[8886] = 8'he4 ;
            rom[8887] = 8'h3b ;
            rom[8888] = 8'hf9 ;
            rom[8889] = 8'h10 ;
            rom[8890] = 8'h18 ;
            rom[8891] = 8'hfd ;
            rom[8892] = 8'h06 ;
            rom[8893] = 8'hca ;
            rom[8894] = 8'he4 ;
            rom[8895] = 8'hd6 ;
            rom[8896] = 8'hea ;
            rom[8897] = 8'he3 ;
            rom[8898] = 8'h36 ;
            rom[8899] = 8'h01 ;
            rom[8900] = 8'hf4 ;
            rom[8901] = 8'hfa ;
            rom[8902] = 8'he9 ;
            rom[8903] = 8'hef ;
            rom[8904] = 8'h0c ;
            rom[8905] = 8'hfe ;
            rom[8906] = 8'h03 ;
            rom[8907] = 8'h46 ;
            rom[8908] = 8'h16 ;
            rom[8909] = 8'hfe ;
            rom[8910] = 8'hfc ;
            rom[8911] = 8'hf7 ;
            rom[8912] = 8'heb ;
            rom[8913] = 8'hf7 ;
            rom[8914] = 8'h15 ;
            rom[8915] = 8'h04 ;
            rom[8916] = 8'hfd ;
            rom[8917] = 8'h0b ;
            rom[8918] = 8'he8 ;
            rom[8919] = 8'hf0 ;
            rom[8920] = 8'h0d ;
            rom[8921] = 8'h0e ;
            rom[8922] = 8'h1b ;
            rom[8923] = 8'h0f ;
            rom[8924] = 8'hfb ;
            rom[8925] = 8'h19 ;
            rom[8926] = 8'h08 ;
            rom[8927] = 8'h0a ;
            rom[8928] = 8'h08 ;
            rom[8929] = 8'h0e ;
            rom[8930] = 8'h29 ;
            rom[8931] = 8'he5 ;
            rom[8932] = 8'h02 ;
            rom[8933] = 8'he8 ;
            rom[8934] = 8'he2 ;
            rom[8935] = 8'hd5 ;
            rom[8936] = 8'hf7 ;
            rom[8937] = 8'hed ;
            rom[8938] = 8'h16 ;
            rom[8939] = 8'h21 ;
            rom[8940] = 8'he3 ;
            rom[8941] = 8'h0f ;
            rom[8942] = 8'hfa ;
            rom[8943] = 8'hef ;
            rom[8944] = 8'hc0 ;
            rom[8945] = 8'h0e ;
            rom[8946] = 8'h16 ;
            rom[8947] = 8'h40 ;
            rom[8948] = 8'hf4 ;
            rom[8949] = 8'hf1 ;
            rom[8950] = 8'h2d ;
            rom[8951] = 8'he2 ;
            rom[8952] = 8'hf0 ;
            rom[8953] = 8'h08 ;
            rom[8954] = 8'hf9 ;
            rom[8955] = 8'h16 ;
            rom[8956] = 8'hf1 ;
            rom[8957] = 8'hd0 ;
            rom[8958] = 8'hfe ;
            rom[8959] = 8'h03 ;
            rom[8960] = 8'h16 ;
            rom[8961] = 8'hde ;
            rom[8962] = 8'hfe ;
            rom[8963] = 8'h02 ;
            rom[8964] = 8'hd3 ;
            rom[8965] = 8'h09 ;
            rom[8966] = 8'hf0 ;
            rom[8967] = 8'h07 ;
            rom[8968] = 8'hf2 ;
            rom[8969] = 8'hf1 ;
            rom[8970] = 8'hed ;
            rom[8971] = 8'h0c ;
            rom[8972] = 8'h1a ;
            rom[8973] = 8'h0b ;
            rom[8974] = 8'h11 ;
            rom[8975] = 8'h00 ;
            rom[8976] = 8'h01 ;
            rom[8977] = 8'hf0 ;
            rom[8978] = 8'h08 ;
            rom[8979] = 8'h22 ;
            rom[8980] = 8'hfd ;
            rom[8981] = 8'hba ;
            rom[8982] = 8'h32 ;
            rom[8983] = 8'heb ;
            rom[8984] = 8'h11 ;
            rom[8985] = 8'hd3 ;
            rom[8986] = 8'h09 ;
            rom[8987] = 8'hcd ;
            rom[8988] = 8'hf9 ;
            rom[8989] = 8'h01 ;
            rom[8990] = 8'hbc ;
            rom[8991] = 8'h0e ;
            rom[8992] = 8'hff ;
            rom[8993] = 8'h0c ;
            rom[8994] = 8'h03 ;
            rom[8995] = 8'he2 ;
            rom[8996] = 8'h07 ;
            rom[8997] = 8'hdd ;
            rom[8998] = 8'hf6 ;
            rom[8999] = 8'hb0 ;
            rom[9000] = 8'h19 ;
            rom[9001] = 8'hdc ;
            rom[9002] = 8'h09 ;
            rom[9003] = 8'hfc ;
            rom[9004] = 8'h0b ;
            rom[9005] = 8'h05 ;
            rom[9006] = 8'hed ;
            rom[9007] = 8'h03 ;
            rom[9008] = 8'he2 ;
            rom[9009] = 8'hfb ;
            rom[9010] = 8'hfb ;
            rom[9011] = 8'hf3 ;
            rom[9012] = 8'hf3 ;
            rom[9013] = 8'hf7 ;
            rom[9014] = 8'hf4 ;
            rom[9015] = 8'h16 ;
            rom[9016] = 8'h0e ;
            rom[9017] = 8'h09 ;
            rom[9018] = 8'hf6 ;
            rom[9019] = 8'he2 ;
            rom[9020] = 8'h15 ;
            rom[9021] = 8'h0d ;
            rom[9022] = 8'hf1 ;
            rom[9023] = 8'he0 ;
            rom[9024] = 8'hf5 ;
            rom[9025] = 8'h0a ;
            rom[9026] = 8'hdb ;
            rom[9027] = 8'hf5 ;
            rom[9028] = 8'h13 ;
            rom[9029] = 8'h18 ;
            rom[9030] = 8'hf5 ;
            rom[9031] = 8'hf6 ;
            rom[9032] = 8'h02 ;
            rom[9033] = 8'hf2 ;
            rom[9034] = 8'he9 ;
            rom[9035] = 8'hfb ;
            rom[9036] = 8'hb3 ;
            rom[9037] = 8'h10 ;
            rom[9038] = 8'h19 ;
            rom[9039] = 8'h12 ;
            rom[9040] = 8'hc3 ;
            rom[9041] = 8'h21 ;
            rom[9042] = 8'hf6 ;
            rom[9043] = 8'he3 ;
            rom[9044] = 8'h16 ;
            rom[9045] = 8'he6 ;
            rom[9046] = 8'he7 ;
            rom[9047] = 8'hf8 ;
            rom[9048] = 8'hc0 ;
            rom[9049] = 8'he2 ;
            rom[9050] = 8'hff ;
            rom[9051] = 8'h00 ;
            rom[9052] = 8'h0c ;
            rom[9053] = 8'hf1 ;
            rom[9054] = 8'h16 ;
            rom[9055] = 8'h00 ;
            rom[9056] = 8'hf9 ;
            rom[9057] = 8'hf5 ;
            rom[9058] = 8'hda ;
            rom[9059] = 8'h25 ;
            rom[9060] = 8'he7 ;
            rom[9061] = 8'h1a ;
            rom[9062] = 8'hfd ;
            rom[9063] = 8'hd4 ;
            rom[9064] = 8'hfe ;
            rom[9065] = 8'h01 ;
            rom[9066] = 8'hf0 ;
            rom[9067] = 8'hfa ;
            rom[9068] = 8'hea ;
            rom[9069] = 8'h06 ;
            rom[9070] = 8'h14 ;
            rom[9071] = 8'he1 ;
            rom[9072] = 8'hfd ;
            rom[9073] = 8'hed ;
            rom[9074] = 8'h12 ;
            rom[9075] = 8'h02 ;
            rom[9076] = 8'hd9 ;
            rom[9077] = 8'h01 ;
            rom[9078] = 8'hf1 ;
            rom[9079] = 8'h03 ;
            rom[9080] = 8'h13 ;
            rom[9081] = 8'hc8 ;
            rom[9082] = 8'hc4 ;
            rom[9083] = 8'h10 ;
            rom[9084] = 8'he6 ;
            rom[9085] = 8'h0a ;
            rom[9086] = 8'hf6 ;
            rom[9087] = 8'h04 ;
            rom[9088] = 8'h0d ;
            rom[9089] = 8'he6 ;
            rom[9090] = 8'he9 ;
            rom[9091] = 8'h06 ;
            rom[9092] = 8'hd4 ;
            rom[9093] = 8'hf5 ;
            rom[9094] = 8'h24 ;
            rom[9095] = 8'hfa ;
            rom[9096] = 8'hdb ;
            rom[9097] = 8'hec ;
            rom[9098] = 8'h26 ;
            rom[9099] = 8'h02 ;
            rom[9100] = 8'hec ;
            rom[9101] = 8'hf5 ;
            rom[9102] = 8'h06 ;
            rom[9103] = 8'he5 ;
            rom[9104] = 8'hfc ;
            rom[9105] = 8'h14 ;
            rom[9106] = 8'h0a ;
            rom[9107] = 8'hfe ;
            rom[9108] = 8'hf4 ;
            rom[9109] = 8'hf5 ;
            rom[9110] = 8'h15 ;
            rom[9111] = 8'hef ;
            rom[9112] = 8'h06 ;
            rom[9113] = 8'he0 ;
            rom[9114] = 8'hf4 ;
            rom[9115] = 8'hc4 ;
            rom[9116] = 8'hfa ;
            rom[9117] = 8'hdb ;
            rom[9118] = 8'h02 ;
            rom[9119] = 8'h0d ;
            rom[9120] = 8'h0e ;
            rom[9121] = 8'h0c ;
            rom[9122] = 8'he4 ;
            rom[9123] = 8'hd7 ;
            rom[9124] = 8'h2a ;
            rom[9125] = 8'he5 ;
            rom[9126] = 8'h0c ;
            rom[9127] = 8'h04 ;
            rom[9128] = 8'h0b ;
            rom[9129] = 8'h05 ;
            rom[9130] = 8'hf3 ;
            rom[9131] = 8'h08 ;
            rom[9132] = 8'h08 ;
            rom[9133] = 8'hfd ;
            rom[9134] = 8'hde ;
            rom[9135] = 8'h1a ;
            rom[9136] = 8'h18 ;
            rom[9137] = 8'h17 ;
            rom[9138] = 8'he5 ;
            rom[9139] = 8'he9 ;
            rom[9140] = 8'he3 ;
            rom[9141] = 8'h0d ;
            rom[9142] = 8'h0e ;
            rom[9143] = 8'h0f ;
            rom[9144] = 8'hdf ;
            rom[9145] = 8'hdb ;
            rom[9146] = 8'hd7 ;
            rom[9147] = 8'h16 ;
            rom[9148] = 8'h40 ;
            rom[9149] = 8'h06 ;
            rom[9150] = 8'hf9 ;
            rom[9151] = 8'hcc ;
            rom[9152] = 8'h0f ;
            rom[9153] = 8'h0c ;
            rom[9154] = 8'h08 ;
            rom[9155] = 8'hf9 ;
            rom[9156] = 8'hff ;
            rom[9157] = 8'h2d ;
            rom[9158] = 8'h00 ;
            rom[9159] = 8'h1b ;
            rom[9160] = 8'he9 ;
            rom[9161] = 8'hfe ;
            rom[9162] = 8'he6 ;
            rom[9163] = 8'hde ;
            rom[9164] = 8'hf7 ;
            rom[9165] = 8'hf6 ;
            rom[9166] = 8'hd9 ;
            rom[9167] = 8'h14 ;
            rom[9168] = 8'h06 ;
            rom[9169] = 8'hd1 ;
            rom[9170] = 8'hf9 ;
            rom[9171] = 8'hed ;
            rom[9172] = 8'hd8 ;
            rom[9173] = 8'hd8 ;
            rom[9174] = 8'h07 ;
            rom[9175] = 8'h25 ;
            rom[9176] = 8'h03 ;
            rom[9177] = 8'h08 ;
            rom[9178] = 8'hf8 ;
            rom[9179] = 8'hff ;
            rom[9180] = 8'ha7 ;
            rom[9181] = 8'h01 ;
            rom[9182] = 8'h05 ;
            rom[9183] = 8'he2 ;
            rom[9184] = 8'h13 ;
            rom[9185] = 8'h3d ;
            rom[9186] = 8'hf1 ;
            rom[9187] = 8'hff ;
            rom[9188] = 8'hcc ;
            rom[9189] = 8'h01 ;
            rom[9190] = 8'h26 ;
            rom[9191] = 8'he0 ;
            rom[9192] = 8'h0a ;
            rom[9193] = 8'h09 ;
            rom[9194] = 8'hf7 ;
            rom[9195] = 8'hdb ;
            rom[9196] = 8'h08 ;
            rom[9197] = 8'h05 ;
            rom[9198] = 8'h04 ;
            rom[9199] = 8'hf2 ;
            rom[9200] = 8'h23 ;
            rom[9201] = 8'h02 ;
            rom[9202] = 8'hf8 ;
            rom[9203] = 8'h01 ;
            rom[9204] = 8'he7 ;
            rom[9205] = 8'h16 ;
            rom[9206] = 8'hff ;
            rom[9207] = 8'h07 ;
            rom[9208] = 8'h06 ;
            rom[9209] = 8'h16 ;
            rom[9210] = 8'hc8 ;
            rom[9211] = 8'hed ;
            rom[9212] = 8'hff ;
            rom[9213] = 8'h2a ;
            rom[9214] = 8'hf1 ;
            rom[9215] = 8'hd8 ;
            rom[9216] = 8'h07 ;
            rom[9217] = 8'hfa ;
            rom[9218] = 8'h2c ;
            rom[9219] = 8'h04 ;
            rom[9220] = 8'hf3 ;
            rom[9221] = 8'he0 ;
            rom[9222] = 8'h0f ;
            rom[9223] = 8'hca ;
            rom[9224] = 8'h2b ;
            rom[9225] = 8'hef ;
            rom[9226] = 8'h0c ;
            rom[9227] = 8'h0f ;
            rom[9228] = 8'h0b ;
            rom[9229] = 8'hec ;
            rom[9230] = 8'he7 ;
            rom[9231] = 8'hda ;
            rom[9232] = 8'hce ;
            rom[9233] = 8'hf5 ;
            rom[9234] = 8'h0c ;
            rom[9235] = 8'hfa ;
            rom[9236] = 8'hf3 ;
            rom[9237] = 8'hdd ;
            rom[9238] = 8'hf6 ;
            rom[9239] = 8'hd4 ;
            rom[9240] = 8'he3 ;
            rom[9241] = 8'hfc ;
            rom[9242] = 8'hf0 ;
            rom[9243] = 8'hbe ;
            rom[9244] = 8'hf9 ;
            rom[9245] = 8'hf0 ;
            rom[9246] = 8'hf5 ;
            rom[9247] = 8'hf8 ;
            rom[9248] = 8'he6 ;
            rom[9249] = 8'hf1 ;
            rom[9250] = 8'hd1 ;
            rom[9251] = 8'hf1 ;
            rom[9252] = 8'he7 ;
            rom[9253] = 8'he9 ;
            rom[9254] = 8'hf8 ;
            rom[9255] = 8'h20 ;
            rom[9256] = 8'hf1 ;
            rom[9257] = 8'h19 ;
            rom[9258] = 8'h0f ;
            rom[9259] = 8'h05 ;
            rom[9260] = 8'hff ;
            rom[9261] = 8'h0c ;
            rom[9262] = 8'hea ;
            rom[9263] = 8'h02 ;
            rom[9264] = 8'he5 ;
            rom[9265] = 8'h04 ;
            rom[9266] = 8'hf9 ;
            rom[9267] = 8'hdb ;
            rom[9268] = 8'h0b ;
            rom[9269] = 8'hed ;
            rom[9270] = 8'hbc ;
            rom[9271] = 8'h12 ;
            rom[9272] = 8'hfc ;
            rom[9273] = 8'h0a ;
            rom[9274] = 8'hd4 ;
            rom[9275] = 8'h04 ;
            rom[9276] = 8'h02 ;
            rom[9277] = 8'h00 ;
            rom[9278] = 8'hf1 ;
            rom[9279] = 8'he7 ;
            rom[9280] = 8'hce ;
            rom[9281] = 8'hfa ;
            rom[9282] = 8'h07 ;
            rom[9283] = 8'h0c ;
            rom[9284] = 8'h09 ;
            rom[9285] = 8'h03 ;
            rom[9286] = 8'hc8 ;
            rom[9287] = 8'h22 ;
            rom[9288] = 8'hfc ;
            rom[9289] = 8'h01 ;
            rom[9290] = 8'hdf ;
            rom[9291] = 8'h0c ;
            rom[9292] = 8'h17 ;
            rom[9293] = 8'hf6 ;
            rom[9294] = 8'he3 ;
            rom[9295] = 8'hcf ;
            rom[9296] = 8'h18 ;
            rom[9297] = 8'hf6 ;
            rom[9298] = 8'hd0 ;
            rom[9299] = 8'h24 ;
            rom[9300] = 8'hef ;
            rom[9301] = 8'hc1 ;
            rom[9302] = 8'hfd ;
            rom[9303] = 8'hfe ;
            rom[9304] = 8'hb5 ;
            rom[9305] = 8'hef ;
            rom[9306] = 8'hdf ;
            rom[9307] = 8'h12 ;
            rom[9308] = 8'hfd ;
            rom[9309] = 8'hd6 ;
            rom[9310] = 8'h10 ;
            rom[9311] = 8'hec ;
            rom[9312] = 8'he0 ;
            rom[9313] = 8'he0 ;
            rom[9314] = 8'hc4 ;
            rom[9315] = 8'h01 ;
            rom[9316] = 8'h0e ;
            rom[9317] = 8'h27 ;
            rom[9318] = 8'hf9 ;
            rom[9319] = 8'ha7 ;
            rom[9320] = 8'hd3 ;
            rom[9321] = 8'h21 ;
            rom[9322] = 8'hed ;
            rom[9323] = 8'h0b ;
            rom[9324] = 8'hdc ;
            rom[9325] = 8'hd9 ;
            rom[9326] = 8'h15 ;
            rom[9327] = 8'hf2 ;
            rom[9328] = 8'hd5 ;
            rom[9329] = 8'hea ;
            rom[9330] = 8'h16 ;
            rom[9331] = 8'hda ;
            rom[9332] = 8'h09 ;
            rom[9333] = 8'h12 ;
            rom[9334] = 8'hd2 ;
            rom[9335] = 8'hf2 ;
            rom[9336] = 8'hf0 ;
            rom[9337] = 8'hbf ;
            rom[9338] = 8'hfb ;
            rom[9339] = 8'h10 ;
            rom[9340] = 8'hdb ;
            rom[9341] = 8'hf7 ;
            rom[9342] = 8'hdc ;
            rom[9343] = 8'he2 ;
            rom[9344] = 8'h03 ;
            rom[9345] = 8'hdd ;
            rom[9346] = 8'hf4 ;
            rom[9347] = 8'h09 ;
            rom[9348] = 8'h17 ;
            rom[9349] = 8'h07 ;
            rom[9350] = 8'hf4 ;
            rom[9351] = 8'hf3 ;
            rom[9352] = 8'hfd ;
            rom[9353] = 8'h20 ;
            rom[9354] = 8'hf3 ;
            rom[9355] = 8'h01 ;
            rom[9356] = 8'hc5 ;
            rom[9357] = 8'hf7 ;
            rom[9358] = 8'h26 ;
            rom[9359] = 8'hef ;
            rom[9360] = 8'h13 ;
            rom[9361] = 8'h04 ;
            rom[9362] = 8'h08 ;
            rom[9363] = 8'h1c ;
            rom[9364] = 8'h16 ;
            rom[9365] = 8'hf1 ;
            rom[9366] = 8'hfd ;
            rom[9367] = 8'hfb ;
            rom[9368] = 8'hc9 ;
            rom[9369] = 8'h07 ;
            rom[9370] = 8'h05 ;
            rom[9371] = 8'hd8 ;
            rom[9372] = 8'hf7 ;
            rom[9373] = 8'hfd ;
            rom[9374] = 8'hde ;
            rom[9375] = 8'hec ;
            rom[9376] = 8'he6 ;
            rom[9377] = 8'h0a ;
            rom[9378] = 8'h13 ;
            rom[9379] = 8'he7 ;
            rom[9380] = 8'h17 ;
            rom[9381] = 8'hf2 ;
            rom[9382] = 8'hf8 ;
            rom[9383] = 8'hc0 ;
            rom[9384] = 8'h09 ;
            rom[9385] = 8'h0f ;
            rom[9386] = 8'hec ;
            rom[9387] = 8'h01 ;
            rom[9388] = 8'h07 ;
            rom[9389] = 8'h1f ;
            rom[9390] = 8'h11 ;
            rom[9391] = 8'hd4 ;
            rom[9392] = 8'he6 ;
            rom[9393] = 8'hc9 ;
            rom[9394] = 8'hff ;
            rom[9395] = 8'hf0 ;
            rom[9396] = 8'h1b ;
            rom[9397] = 8'hd8 ;
            rom[9398] = 8'he8 ;
            rom[9399] = 8'h0f ;
            rom[9400] = 8'h22 ;
            rom[9401] = 8'hf9 ;
            rom[9402] = 8'h0c ;
            rom[9403] = 8'hed ;
            rom[9404] = 8'hfe ;
            rom[9405] = 8'hd3 ;
            rom[9406] = 8'h00 ;
            rom[9407] = 8'h07 ;
            rom[9408] = 8'hf1 ;
            rom[9409] = 8'hf2 ;
            rom[9410] = 8'hfa ;
            rom[9411] = 8'hc3 ;
            rom[9412] = 8'hd7 ;
            rom[9413] = 8'hdf ;
            rom[9414] = 8'hef ;
            rom[9415] = 8'h01 ;
            rom[9416] = 8'hea ;
            rom[9417] = 8'h04 ;
            rom[9418] = 8'hff ;
            rom[9419] = 8'h08 ;
            rom[9420] = 8'he1 ;
            rom[9421] = 8'h25 ;
            rom[9422] = 8'hef ;
            rom[9423] = 8'h10 ;
            rom[9424] = 8'hdc ;
            rom[9425] = 8'h30 ;
            rom[9426] = 8'hfc ;
            rom[9427] = 8'hf3 ;
            rom[9428] = 8'h13 ;
            rom[9429] = 8'h1d ;
            rom[9430] = 8'h08 ;
            rom[9431] = 8'he2 ;
            rom[9432] = 8'h21 ;
            rom[9433] = 8'heb ;
            rom[9434] = 8'h06 ;
            rom[9435] = 8'hee ;
            rom[9436] = 8'hce ;
            rom[9437] = 8'h04 ;
            rom[9438] = 8'h04 ;
            rom[9439] = 8'h21 ;
            rom[9440] = 8'hf8 ;
            rom[9441] = 8'h11 ;
            rom[9442] = 8'h10 ;
            rom[9443] = 8'h01 ;
            rom[9444] = 8'hed ;
            rom[9445] = 8'hc8 ;
            rom[9446] = 8'hc8 ;
            rom[9447] = 8'h02 ;
            rom[9448] = 8'h01 ;
            rom[9449] = 8'hf5 ;
            rom[9450] = 8'he8 ;
            rom[9451] = 8'hf0 ;
            rom[9452] = 8'he4 ;
            rom[9453] = 8'hd8 ;
            rom[9454] = 8'h0e ;
            rom[9455] = 8'he5 ;
            rom[9456] = 8'hef ;
            rom[9457] = 8'h0c ;
            rom[9458] = 8'h0e ;
            rom[9459] = 8'hfa ;
            rom[9460] = 8'h00 ;
            rom[9461] = 8'h29 ;
            rom[9462] = 8'h15 ;
            rom[9463] = 8'h0d ;
            rom[9464] = 8'h11 ;
            rom[9465] = 8'h0f ;
            rom[9466] = 8'h12 ;
            rom[9467] = 8'h0e ;
            rom[9468] = 8'hf8 ;
            rom[9469] = 8'he6 ;
            rom[9470] = 8'he0 ;
            rom[9471] = 8'hc8 ;
            rom[9472] = 8'hd7 ;
            rom[9473] = 8'h03 ;
            rom[9474] = 8'he6 ;
            rom[9475] = 8'h14 ;
            rom[9476] = 8'hf5 ;
            rom[9477] = 8'hfb ;
            rom[9478] = 8'he7 ;
            rom[9479] = 8'hd5 ;
            rom[9480] = 8'h12 ;
            rom[9481] = 8'hfb ;
            rom[9482] = 8'h14 ;
            rom[9483] = 8'hf4 ;
            rom[9484] = 8'hf1 ;
            rom[9485] = 8'he8 ;
            rom[9486] = 8'h1f ;
            rom[9487] = 8'h00 ;
            rom[9488] = 8'hec ;
            rom[9489] = 8'h05 ;
            rom[9490] = 8'he8 ;
            rom[9491] = 8'hf0 ;
            rom[9492] = 8'hf4 ;
            rom[9493] = 8'h15 ;
            rom[9494] = 8'h0a ;
            rom[9495] = 8'hf2 ;
            rom[9496] = 8'h0c ;
            rom[9497] = 8'hee ;
            rom[9498] = 8'h08 ;
            rom[9499] = 8'h08 ;
            rom[9500] = 8'he2 ;
            rom[9501] = 8'h0b ;
            rom[9502] = 8'h34 ;
            rom[9503] = 8'h05 ;
            rom[9504] = 8'h0b ;
            rom[9505] = 8'hed ;
            rom[9506] = 8'hc7 ;
            rom[9507] = 8'hd8 ;
            rom[9508] = 8'hfd ;
            rom[9509] = 8'hec ;
            rom[9510] = 8'hf7 ;
            rom[9511] = 8'h04 ;
            rom[9512] = 8'hf5 ;
            rom[9513] = 8'heb ;
            rom[9514] = 8'h03 ;
            rom[9515] = 8'h1c ;
            rom[9516] = 8'h22 ;
            rom[9517] = 8'hea ;
            rom[9518] = 8'h08 ;
            rom[9519] = 8'hc5 ;
            rom[9520] = 8'hed ;
            rom[9521] = 8'h32 ;
            rom[9522] = 8'h00 ;
            rom[9523] = 8'hf2 ;
            rom[9524] = 8'hfb ;
            rom[9525] = 8'h03 ;
            rom[9526] = 8'h0c ;
            rom[9527] = 8'heb ;
            rom[9528] = 8'h1c ;
            rom[9529] = 8'h0d ;
            rom[9530] = 8'h1c ;
            rom[9531] = 8'h15 ;
            rom[9532] = 8'he9 ;
            rom[9533] = 8'hdd ;
            rom[9534] = 8'h06 ;
            rom[9535] = 8'h02 ;
            rom[9536] = 8'h07 ;
            rom[9537] = 8'h15 ;
            rom[9538] = 8'h0e ;
            rom[9539] = 8'hd5 ;
            rom[9540] = 8'h12 ;
            rom[9541] = 8'he9 ;
            rom[9542] = 8'he0 ;
            rom[9543] = 8'hf8 ;
            rom[9544] = 8'h04 ;
            rom[9545] = 8'he9 ;
            rom[9546] = 8'hd1 ;
            rom[9547] = 8'hf9 ;
            rom[9548] = 8'hc4 ;
            rom[9549] = 8'h07 ;
            rom[9550] = 8'hdf ;
            rom[9551] = 8'h01 ;
            rom[9552] = 8'h25 ;
            rom[9553] = 8'h28 ;
            rom[9554] = 8'h0a ;
            rom[9555] = 8'hf2 ;
            rom[9556] = 8'h02 ;
            rom[9557] = 8'heb ;
            rom[9558] = 8'hd5 ;
            rom[9559] = 8'he0 ;
            rom[9560] = 8'hf7 ;
            rom[9561] = 8'h31 ;
            rom[9562] = 8'hd6 ;
            rom[9563] = 8'h02 ;
            rom[9564] = 8'he7 ;
            rom[9565] = 8'hfb ;
            rom[9566] = 8'hcf ;
            rom[9567] = 8'hc1 ;
            rom[9568] = 8'h03 ;
            rom[9569] = 8'h0e ;
            rom[9570] = 8'h01 ;
            rom[9571] = 8'he8 ;
            rom[9572] = 8'h05 ;
            rom[9573] = 8'hfd ;
            rom[9574] = 8'h0b ;
            rom[9575] = 8'h18 ;
            rom[9576] = 8'he8 ;
            rom[9577] = 8'h0b ;
            rom[9578] = 8'h00 ;
            rom[9579] = 8'h09 ;
            rom[9580] = 8'hfc ;
            rom[9581] = 8'he7 ;
            rom[9582] = 8'hda ;
            rom[9583] = 8'h05 ;
            rom[9584] = 8'h16 ;
            rom[9585] = 8'he8 ;
            rom[9586] = 8'h11 ;
            rom[9587] = 8'hfc ;
            rom[9588] = 8'h27 ;
            rom[9589] = 8'h11 ;
            rom[9590] = 8'h20 ;
            rom[9591] = 8'h00 ;
            rom[9592] = 8'h0c ;
            rom[9593] = 8'h2d ;
            rom[9594] = 8'hfa ;
            rom[9595] = 8'hdd ;
            rom[9596] = 8'hfa ;
            rom[9597] = 8'hf8 ;
            rom[9598] = 8'h00 ;
            rom[9599] = 8'h04 ;
            rom[9600] = 8'hd9 ;
            rom[9601] = 8'h00 ;
            rom[9602] = 8'he1 ;
            rom[9603] = 8'hf8 ;
            rom[9604] = 8'hdb ;
            rom[9605] = 8'hf0 ;
            rom[9606] = 8'h01 ;
            rom[9607] = 8'hfe ;
            rom[9608] = 8'hf4 ;
            rom[9609] = 8'hf8 ;
            rom[9610] = 8'h0c ;
            rom[9611] = 8'hce ;
            rom[9612] = 8'hfd ;
            rom[9613] = 8'h09 ;
            rom[9614] = 8'h08 ;
            rom[9615] = 8'hc7 ;
            rom[9616] = 8'hfc ;
            rom[9617] = 8'hf8 ;
            rom[9618] = 8'hfd ;
            rom[9619] = 8'he8 ;
            rom[9620] = 8'hf4 ;
            rom[9621] = 8'hfe ;
            rom[9622] = 8'h0e ;
            rom[9623] = 8'hec ;
            rom[9624] = 8'h0d ;
            rom[9625] = 8'h03 ;
            rom[9626] = 8'hb3 ;
            rom[9627] = 8'h00 ;
            rom[9628] = 8'h11 ;
            rom[9629] = 8'hf7 ;
            rom[9630] = 8'h0f ;
            rom[9631] = 8'heb ;
            rom[9632] = 8'hfe ;
            rom[9633] = 8'h13 ;
            rom[9634] = 8'hec ;
            rom[9635] = 8'h00 ;
            rom[9636] = 8'hf3 ;
            rom[9637] = 8'heb ;
            rom[9638] = 8'h23 ;
            rom[9639] = 8'hec ;
            rom[9640] = 8'hc2 ;
            rom[9641] = 8'hd6 ;
            rom[9642] = 8'he3 ;
            rom[9643] = 8'h05 ;
            rom[9644] = 8'h1f ;
            rom[9645] = 8'hd3 ;
            rom[9646] = 8'h02 ;
            rom[9647] = 8'he4 ;
            rom[9648] = 8'h13 ;
            rom[9649] = 8'h0c ;
            rom[9650] = 8'hbe ;
            rom[9651] = 8'he9 ;
            rom[9652] = 8'he4 ;
            rom[9653] = 8'hf5 ;
            rom[9654] = 8'h04 ;
            rom[9655] = 8'h05 ;
            rom[9656] = 8'h0a ;
            rom[9657] = 8'hf4 ;
            rom[9658] = 8'h0b ;
            rom[9659] = 8'hea ;
            rom[9660] = 8'hfa ;
            rom[9661] = 8'hf0 ;
            rom[9662] = 8'hf7 ;
            rom[9663] = 8'he9 ;
            rom[9664] = 8'h14 ;
            rom[9665] = 8'h06 ;
            rom[9666] = 8'hf7 ;
            rom[9667] = 8'hc7 ;
            rom[9668] = 8'hf7 ;
            rom[9669] = 8'hf4 ;
            rom[9670] = 8'hf3 ;
            rom[9671] = 8'hc8 ;
            rom[9672] = 8'he0 ;
            rom[9673] = 8'hef ;
            rom[9674] = 8'hb5 ;
            rom[9675] = 8'hf5 ;
            rom[9676] = 8'hee ;
            rom[9677] = 8'hff ;
            rom[9678] = 8'he6 ;
            rom[9679] = 8'h11 ;
            rom[9680] = 8'h12 ;
            rom[9681] = 8'h04 ;
            rom[9682] = 8'hf5 ;
            rom[9683] = 8'hf9 ;
            rom[9684] = 8'hfe ;
            rom[9685] = 8'hf0 ;
            rom[9686] = 8'hf5 ;
            rom[9687] = 8'h00 ;
            rom[9688] = 8'h06 ;
            rom[9689] = 8'h0e ;
            rom[9690] = 8'hf7 ;
            rom[9691] = 8'h21 ;
            rom[9692] = 8'he2 ;
            rom[9693] = 8'h02 ;
            rom[9694] = 8'hd8 ;
            rom[9695] = 8'hef ;
            rom[9696] = 8'h06 ;
            rom[9697] = 8'h02 ;
            rom[9698] = 8'hfb ;
            rom[9699] = 8'h07 ;
            rom[9700] = 8'h13 ;
            rom[9701] = 8'hfa ;
            rom[9702] = 8'hfb ;
            rom[9703] = 8'h15 ;
            rom[9704] = 8'he4 ;
            rom[9705] = 8'h07 ;
            rom[9706] = 8'hfc ;
            rom[9707] = 8'hfb ;
            rom[9708] = 8'h0f ;
            rom[9709] = 8'h04 ;
            rom[9710] = 8'hea ;
            rom[9711] = 8'h00 ;
            rom[9712] = 8'h09 ;
            rom[9713] = 8'hdd ;
            rom[9714] = 8'h0e ;
            rom[9715] = 8'he0 ;
            rom[9716] = 8'h16 ;
            rom[9717] = 8'h02 ;
            rom[9718] = 8'hca ;
            rom[9719] = 8'hf4 ;
            rom[9720] = 8'he9 ;
            rom[9721] = 8'hf9 ;
            rom[9722] = 8'h02 ;
            rom[9723] = 8'h04 ;
            rom[9724] = 8'h03 ;
            rom[9725] = 8'hf9 ;
            rom[9726] = 8'hff ;
            rom[9727] = 8'hee ;
            rom[9728] = 8'hd8 ;
            rom[9729] = 8'hf8 ;
            rom[9730] = 8'h0f ;
            rom[9731] = 8'hda ;
            rom[9732] = 8'he0 ;
            rom[9733] = 8'h24 ;
            rom[9734] = 8'he7 ;
            rom[9735] = 8'h12 ;
            rom[9736] = 8'hfb ;
            rom[9737] = 8'he8 ;
            rom[9738] = 8'hf9 ;
            rom[9739] = 8'hf4 ;
            rom[9740] = 8'h42 ;
            rom[9741] = 8'h09 ;
            rom[9742] = 8'h32 ;
            rom[9743] = 8'h00 ;
            rom[9744] = 8'h12 ;
            rom[9745] = 8'heb ;
            rom[9746] = 8'hf2 ;
            rom[9747] = 8'h15 ;
            rom[9748] = 8'he1 ;
            rom[9749] = 8'h01 ;
            rom[9750] = 8'h1d ;
            rom[9751] = 8'hf4 ;
            rom[9752] = 8'h33 ;
            rom[9753] = 8'hf8 ;
            rom[9754] = 8'h17 ;
            rom[9755] = 8'h19 ;
            rom[9756] = 8'hf0 ;
            rom[9757] = 8'h1e ;
            rom[9758] = 8'hf7 ;
            rom[9759] = 8'hd8 ;
            rom[9760] = 8'h07 ;
            rom[9761] = 8'hdf ;
            rom[9762] = 8'hfd ;
            rom[9763] = 8'he8 ;
            rom[9764] = 8'h06 ;
            rom[9765] = 8'h01 ;
            rom[9766] = 8'h05 ;
            rom[9767] = 8'hdf ;
            rom[9768] = 8'h17 ;
            rom[9769] = 8'he2 ;
            rom[9770] = 8'h09 ;
            rom[9771] = 8'h01 ;
            rom[9772] = 8'h00 ;
            rom[9773] = 8'hf8 ;
            rom[9774] = 8'hc7 ;
            rom[9775] = 8'hd6 ;
            rom[9776] = 8'h12 ;
            rom[9777] = 8'h23 ;
            rom[9778] = 8'h2c ;
            rom[9779] = 8'heb ;
            rom[9780] = 8'he5 ;
            rom[9781] = 8'hee ;
            rom[9782] = 8'h25 ;
            rom[9783] = 8'hed ;
            rom[9784] = 8'h05 ;
            rom[9785] = 8'h07 ;
            rom[9786] = 8'h11 ;
            rom[9787] = 8'hf0 ;
            rom[9788] = 8'h01 ;
            rom[9789] = 8'hf3 ;
            rom[9790] = 8'h0d ;
            rom[9791] = 8'h02 ;
            rom[9792] = 8'h05 ;
            rom[9793] = 8'hd0 ;
            rom[9794] = 8'hfe ;
            rom[9795] = 8'h09 ;
            rom[9796] = 8'he7 ;
            rom[9797] = 8'h0a ;
            rom[9798] = 8'h1e ;
            rom[9799] = 8'h03 ;
            rom[9800] = 8'he5 ;
            rom[9801] = 8'hfa ;
            rom[9802] = 8'h00 ;
            rom[9803] = 8'h08 ;
            rom[9804] = 8'hfa ;
            rom[9805] = 8'h02 ;
            rom[9806] = 8'hfb ;
            rom[9807] = 8'hdb ;
            rom[9808] = 8'h14 ;
            rom[9809] = 8'h0c ;
            rom[9810] = 8'hf2 ;
            rom[9811] = 8'he5 ;
            rom[9812] = 8'hfd ;
            rom[9813] = 8'h0e ;
            rom[9814] = 8'hf0 ;
            rom[9815] = 8'hec ;
            rom[9816] = 8'hf1 ;
            rom[9817] = 8'h0d ;
            rom[9818] = 8'he8 ;
            rom[9819] = 8'h0c ;
            rom[9820] = 8'h12 ;
            rom[9821] = 8'hf5 ;
            rom[9822] = 8'hf3 ;
            rom[9823] = 8'hdc ;
            rom[9824] = 8'h18 ;
            rom[9825] = 8'h0f ;
            rom[9826] = 8'hc5 ;
            rom[9827] = 8'h13 ;
            rom[9828] = 8'h20 ;
            rom[9829] = 8'h01 ;
            rom[9830] = 8'hfa ;
            rom[9831] = 8'h10 ;
            rom[9832] = 8'h09 ;
            rom[9833] = 8'h1c ;
            rom[9834] = 8'hea ;
            rom[9835] = 8'h00 ;
            rom[9836] = 8'h14 ;
            rom[9837] = 8'h2a ;
            rom[9838] = 8'hc9 ;
            rom[9839] = 8'h1a ;
            rom[9840] = 8'h15 ;
            rom[9841] = 8'hf1 ;
            rom[9842] = 8'h0d ;
            rom[9843] = 8'he2 ;
            rom[9844] = 8'hf1 ;
            rom[9845] = 8'h05 ;
            rom[9846] = 8'he5 ;
            rom[9847] = 8'h06 ;
            rom[9848] = 8'hfb ;
            rom[9849] = 8'hea ;
            rom[9850] = 8'h0d ;
            rom[9851] = 8'hd4 ;
            rom[9852] = 8'hf3 ;
            rom[9853] = 8'heb ;
            rom[9854] = 8'hff ;
            rom[9855] = 8'h18 ;
            rom[9856] = 8'hec ;
            rom[9857] = 8'hf4 ;
            rom[9858] = 8'hf8 ;
            rom[9859] = 8'h08 ;
            rom[9860] = 8'h13 ;
            rom[9861] = 8'h03 ;
            rom[9862] = 8'hef ;
            rom[9863] = 8'hfd ;
            rom[9864] = 8'h31 ;
            rom[9865] = 8'hdd ;
            rom[9866] = 8'h0b ;
            rom[9867] = 8'hf6 ;
            rom[9868] = 8'hfc ;
            rom[9869] = 8'hdf ;
            rom[9870] = 8'h0a ;
            rom[9871] = 8'hf5 ;
            rom[9872] = 8'hfd ;
            rom[9873] = 8'h0f ;
            rom[9874] = 8'h09 ;
            rom[9875] = 8'h0c ;
            rom[9876] = 8'he7 ;
            rom[9877] = 8'h16 ;
            rom[9878] = 8'he4 ;
            rom[9879] = 8'h00 ;
            rom[9880] = 8'h16 ;
            rom[9881] = 8'h09 ;
            rom[9882] = 8'h14 ;
            rom[9883] = 8'hf9 ;
            rom[9884] = 8'hfd ;
            rom[9885] = 8'h11 ;
            rom[9886] = 8'h00 ;
            rom[9887] = 8'h06 ;
            rom[9888] = 8'h22 ;
            rom[9889] = 8'h16 ;
            rom[9890] = 8'he8 ;
            rom[9891] = 8'hdf ;
            rom[9892] = 8'hc9 ;
            rom[9893] = 8'h07 ;
            rom[9894] = 8'hf5 ;
            rom[9895] = 8'h07 ;
            rom[9896] = 8'h0e ;
            rom[9897] = 8'h08 ;
            rom[9898] = 8'he6 ;
            rom[9899] = 8'hdf ;
            rom[9900] = 8'h26 ;
            rom[9901] = 8'he1 ;
            rom[9902] = 8'hfa ;
            rom[9903] = 8'he9 ;
            rom[9904] = 8'hd6 ;
            rom[9905] = 8'h14 ;
            rom[9906] = 8'he3 ;
            rom[9907] = 8'he1 ;
            rom[9908] = 8'hf4 ;
            rom[9909] = 8'h14 ;
            rom[9910] = 8'h13 ;
            rom[9911] = 8'h15 ;
            rom[9912] = 8'h00 ;
            rom[9913] = 8'h0c ;
            rom[9914] = 8'hef ;
            rom[9915] = 8'hee ;
            rom[9916] = 8'hf9 ;
            rom[9917] = 8'hf7 ;
            rom[9918] = 8'hfe ;
            rom[9919] = 8'he7 ;
            rom[9920] = 8'h26 ;
            rom[9921] = 8'he4 ;
            rom[9922] = 8'h0f ;
            rom[9923] = 8'hf5 ;
            rom[9924] = 8'hf4 ;
            rom[9925] = 8'hf6 ;
            rom[9926] = 8'heb ;
            rom[9927] = 8'he8 ;
            rom[9928] = 8'h03 ;
            rom[9929] = 8'hfa ;
            rom[9930] = 8'heb ;
            rom[9931] = 8'he3 ;
            rom[9932] = 8'h0c ;
            rom[9933] = 8'hdf ;
            rom[9934] = 8'h00 ;
            rom[9935] = 8'h0b ;
            rom[9936] = 8'heb ;
            rom[9937] = 8'h0a ;
            rom[9938] = 8'hef ;
            rom[9939] = 8'heb ;
            rom[9940] = 8'hfa ;
            rom[9941] = 8'he5 ;
            rom[9942] = 8'hfe ;
            rom[9943] = 8'hcf ;
            rom[9944] = 8'hfe ;
            rom[9945] = 8'h09 ;
            rom[9946] = 8'hfa ;
            rom[9947] = 8'h05 ;
            rom[9948] = 8'hf5 ;
            rom[9949] = 8'h0f ;
            rom[9950] = 8'h02 ;
            rom[9951] = 8'hf8 ;
            rom[9952] = 8'h0f ;
            rom[9953] = 8'h07 ;
            rom[9954] = 8'h06 ;
            rom[9955] = 8'hd8 ;
            rom[9956] = 8'h08 ;
            rom[9957] = 8'hbe ;
            rom[9958] = 8'h0c ;
            rom[9959] = 8'hf5 ;
            rom[9960] = 8'h35 ;
            rom[9961] = 8'h24 ;
            rom[9962] = 8'h06 ;
            rom[9963] = 8'h12 ;
            rom[9964] = 8'h0f ;
            rom[9965] = 8'h06 ;
            rom[9966] = 8'h01 ;
            rom[9967] = 8'h05 ;
            rom[9968] = 8'he3 ;
            rom[9969] = 8'he7 ;
            rom[9970] = 8'hfb ;
            rom[9971] = 8'hf5 ;
            rom[9972] = 8'h35 ;
            rom[9973] = 8'hef ;
            rom[9974] = 8'h02 ;
            rom[9975] = 8'h14 ;
            rom[9976] = 8'he9 ;
            rom[9977] = 8'h01 ;
            rom[9978] = 8'h1a ;
            rom[9979] = 8'h03 ;
            rom[9980] = 8'he1 ;
            rom[9981] = 8'h29 ;
            rom[9982] = 8'h1a ;
            rom[9983] = 8'he4 ;
            rom[9984] = 8'hea ;
            rom[9985] = 8'he7 ;
            rom[9986] = 8'hfb ;
            rom[9987] = 8'h20 ;
            rom[9988] = 8'h05 ;
            rom[9989] = 8'hd7 ;
            rom[9990] = 8'h00 ;
            rom[9991] = 8'hd4 ;
            rom[9992] = 8'h2d ;
            rom[9993] = 8'h1d ;
            rom[9994] = 8'hda ;
            rom[9995] = 8'hb2 ;
            rom[9996] = 8'hda ;
            rom[9997] = 8'h08 ;
            rom[9998] = 8'hf1 ;
            rom[9999] = 8'hf4 ;
            rom[10000] = 8'hff ;
            rom[10001] = 8'h02 ;
            rom[10002] = 8'hf2 ;
            rom[10003] = 8'he2 ;
            rom[10004] = 8'hee ;
            rom[10005] = 8'hf0 ;
            rom[10006] = 8'hf6 ;
            rom[10007] = 8'h03 ;
            rom[10008] = 8'h00 ;
            rom[10009] = 8'h09 ;
            rom[10010] = 8'h07 ;
            rom[10011] = 8'h1d ;
            rom[10012] = 8'hf0 ;
            rom[10013] = 8'hf7 ;
            rom[10014] = 8'h05 ;
            rom[10015] = 8'hbe ;
            rom[10016] = 8'hd3 ;
            rom[10017] = 8'h09 ;
            rom[10018] = 8'hd4 ;
            rom[10019] = 8'h0b ;
            rom[10020] = 8'hc3 ;
            rom[10021] = 8'h1f ;
            rom[10022] = 8'h16 ;
            rom[10023] = 8'h20 ;
            rom[10024] = 8'hd5 ;
            rom[10025] = 8'he5 ;
            rom[10026] = 8'hf3 ;
            rom[10027] = 8'hd8 ;
            rom[10028] = 8'h37 ;
            rom[10029] = 8'h09 ;
            rom[10030] = 8'h09 ;
            rom[10031] = 8'he1 ;
            rom[10032] = 8'hf7 ;
            rom[10033] = 8'hf9 ;
            rom[10034] = 8'h0a ;
            rom[10035] = 8'hd9 ;
            rom[10036] = 8'h22 ;
            rom[10037] = 8'hf7 ;
            rom[10038] = 8'hdc ;
            rom[10039] = 8'heb ;
            rom[10040] = 8'h07 ;
            rom[10041] = 8'h00 ;
            rom[10042] = 8'h04 ;
            rom[10043] = 8'hd4 ;
            rom[10044] = 8'he9 ;
            rom[10045] = 8'h0d ;
            rom[10046] = 8'he0 ;
            rom[10047] = 8'hf3 ;
            rom[10048] = 8'he1 ;
            rom[10049] = 8'hf0 ;
            rom[10050] = 8'h08 ;
            rom[10051] = 8'heb ;
            rom[10052] = 8'h05 ;
            rom[10053] = 8'he0 ;
            rom[10054] = 8'hdc ;
            rom[10055] = 8'hc8 ;
            rom[10056] = 8'hfe ;
            rom[10057] = 8'he5 ;
            rom[10058] = 8'hf0 ;
            rom[10059] = 8'h1e ;
            rom[10060] = 8'h0c ;
            rom[10061] = 8'he1 ;
            rom[10062] = 8'h1d ;
            rom[10063] = 8'hf9 ;
            rom[10064] = 8'h04 ;
            rom[10065] = 8'he6 ;
            rom[10066] = 8'h07 ;
            rom[10067] = 8'hfc ;
            rom[10068] = 8'h00 ;
            rom[10069] = 8'hed ;
            rom[10070] = 8'he8 ;
            rom[10071] = 8'hfa ;
            rom[10072] = 8'h30 ;
            rom[10073] = 8'h07 ;
            rom[10074] = 8'h0b ;
            rom[10075] = 8'h0f ;
            rom[10076] = 8'h09 ;
            rom[10077] = 8'h07 ;
            rom[10078] = 8'hf9 ;
            rom[10079] = 8'h00 ;
            rom[10080] = 8'hed ;
            rom[10081] = 8'he6 ;
            rom[10082] = 8'h0d ;
            rom[10083] = 8'he8 ;
            rom[10084] = 8'h17 ;
            rom[10085] = 8'hf4 ;
            rom[10086] = 8'h0a ;
            rom[10087] = 8'hfd ;
            rom[10088] = 8'hec ;
            rom[10089] = 8'hb9 ;
            rom[10090] = 8'h04 ;
            rom[10091] = 8'hea ;
            rom[10092] = 8'hf9 ;
            rom[10093] = 8'h1b ;
            rom[10094] = 8'hf6 ;
            rom[10095] = 8'hf8 ;
            rom[10096] = 8'h10 ;
            rom[10097] = 8'hed ;
            rom[10098] = 8'h20 ;
            rom[10099] = 8'h10 ;
            rom[10100] = 8'h0c ;
            rom[10101] = 8'h06 ;
            rom[10102] = 8'h1e ;
            rom[10103] = 8'hf6 ;
            rom[10104] = 8'hf9 ;
            rom[10105] = 8'hfc ;
            rom[10106] = 8'h13 ;
            rom[10107] = 8'h18 ;
            rom[10108] = 8'hf2 ;
            rom[10109] = 8'he6 ;
            rom[10110] = 8'hf2 ;
            rom[10111] = 8'h07 ;
            rom[10112] = 8'hd6 ;
            rom[10113] = 8'he7 ;
            rom[10114] = 8'h07 ;
            rom[10115] = 8'h27 ;
            rom[10116] = 8'h06 ;
            rom[10117] = 8'he3 ;
            rom[10118] = 8'h20 ;
            rom[10119] = 8'hf5 ;
            rom[10120] = 8'hd3 ;
            rom[10121] = 8'hd8 ;
            rom[10122] = 8'hde ;
            rom[10123] = 8'hf4 ;
            rom[10124] = 8'hfb ;
            rom[10125] = 8'h2a ;
            rom[10126] = 8'hf5 ;
            rom[10127] = 8'h00 ;
            rom[10128] = 8'he8 ;
            rom[10129] = 8'hef ;
            rom[10130] = 8'hf1 ;
            rom[10131] = 8'hd7 ;
            rom[10132] = 8'h1d ;
            rom[10133] = 8'hf7 ;
            rom[10134] = 8'hdd ;
            rom[10135] = 8'h12 ;
            rom[10136] = 8'h15 ;
            rom[10137] = 8'hf0 ;
            rom[10138] = 8'hfb ;
            rom[10139] = 8'hec ;
            rom[10140] = 8'h0d ;
            rom[10141] = 8'hec ;
            rom[10142] = 8'h2a ;
            rom[10143] = 8'h0c ;
            rom[10144] = 8'h18 ;
            rom[10145] = 8'hfa ;
            rom[10146] = 8'hfc ;
            rom[10147] = 8'hf0 ;
            rom[10148] = 8'hfb ;
            rom[10149] = 8'h11 ;
            rom[10150] = 8'hf6 ;
            rom[10151] = 8'hf1 ;
            rom[10152] = 8'h08 ;
            rom[10153] = 8'hf8 ;
            rom[10154] = 8'hf7 ;
            rom[10155] = 8'h0b ;
            rom[10156] = 8'h13 ;
            rom[10157] = 8'h08 ;
            rom[10158] = 8'hdd ;
            rom[10159] = 8'h10 ;
            rom[10160] = 8'h1b ;
            rom[10161] = 8'hf9 ;
            rom[10162] = 8'hfe ;
            rom[10163] = 8'h1c ;
            rom[10164] = 8'hf2 ;
            rom[10165] = 8'hf1 ;
            rom[10166] = 8'h08 ;
            rom[10167] = 8'he8 ;
            rom[10168] = 8'hee ;
            rom[10169] = 8'hea ;
            rom[10170] = 8'hfb ;
            rom[10171] = 8'h18 ;
            rom[10172] = 8'h06 ;
            rom[10173] = 8'hf9 ;
            rom[10174] = 8'he5 ;
            rom[10175] = 8'he9 ;
            rom[10176] = 8'hea ;
            rom[10177] = 8'h18 ;
            rom[10178] = 8'he6 ;
            rom[10179] = 8'hed ;
            rom[10180] = 8'h16 ;
            rom[10181] = 8'he6 ;
            rom[10182] = 8'h14 ;
            rom[10183] = 8'h12 ;
            rom[10184] = 8'hfe ;
            rom[10185] = 8'he1 ;
            rom[10186] = 8'h10 ;
            rom[10187] = 8'h11 ;
            rom[10188] = 8'h12 ;
            rom[10189] = 8'hcb ;
            rom[10190] = 8'he9 ;
            rom[10191] = 8'he8 ;
            rom[10192] = 8'h1e ;
            rom[10193] = 8'h03 ;
            rom[10194] = 8'h08 ;
            rom[10195] = 8'hff ;
            rom[10196] = 8'hee ;
            rom[10197] = 8'h14 ;
            rom[10198] = 8'h08 ;
            rom[10199] = 8'heb ;
            rom[10200] = 8'h2e ;
            rom[10201] = 8'hfc ;
            rom[10202] = 8'h12 ;
            rom[10203] = 8'h14 ;
            rom[10204] = 8'hf6 ;
            rom[10205] = 8'h36 ;
            rom[10206] = 8'hf2 ;
            rom[10207] = 8'hfe ;
            rom[10208] = 8'he6 ;
            rom[10209] = 8'h2b ;
            rom[10210] = 8'he8 ;
            rom[10211] = 8'he3 ;
            rom[10212] = 8'h06 ;
            rom[10213] = 8'h0c ;
            rom[10214] = 8'h2f ;
            rom[10215] = 8'hd9 ;
            rom[10216] = 8'hf8 ;
            rom[10217] = 8'hf8 ;
            rom[10218] = 8'h15 ;
            rom[10219] = 8'hf1 ;
            rom[10220] = 8'he3 ;
            rom[10221] = 8'h03 ;
            rom[10222] = 8'hc3 ;
            rom[10223] = 8'h24 ;
            rom[10224] = 8'h10 ;
            rom[10225] = 8'hf8 ;
            rom[10226] = 8'hfa ;
            rom[10227] = 8'h09 ;
            rom[10228] = 8'hfb ;
            rom[10229] = 8'h05 ;
            rom[10230] = 8'h0a ;
            rom[10231] = 8'hf6 ;
            rom[10232] = 8'hef ;
            rom[10233] = 8'h19 ;
            rom[10234] = 8'hfc ;
            rom[10235] = 8'hf8 ;
            rom[10236] = 8'h24 ;
            rom[10237] = 8'h25 ;
            rom[10238] = 8'hfd ;
            rom[10239] = 8'hf4 ;
            rom[10240] = 8'he1 ;
            rom[10241] = 8'heb ;
            rom[10242] = 8'hdb ;
            rom[10243] = 8'h18 ;
            rom[10244] = 8'hfc ;
            rom[10245] = 8'h12 ;
            rom[10246] = 8'h06 ;
            rom[10247] = 8'h05 ;
            rom[10248] = 8'h16 ;
            rom[10249] = 8'hf9 ;
            rom[10250] = 8'hf0 ;
            rom[10251] = 8'hdd ;
            rom[10252] = 8'hef ;
            rom[10253] = 8'hea ;
            rom[10254] = 8'h07 ;
            rom[10255] = 8'h06 ;
            rom[10256] = 8'h07 ;
            rom[10257] = 8'h18 ;
            rom[10258] = 8'hf9 ;
            rom[10259] = 8'hf3 ;
            rom[10260] = 8'h10 ;
            rom[10261] = 8'h0c ;
            rom[10262] = 8'he8 ;
            rom[10263] = 8'h0c ;
            rom[10264] = 8'hef ;
            rom[10265] = 8'hde ;
            rom[10266] = 8'h03 ;
            rom[10267] = 8'hf3 ;
            rom[10268] = 8'hfc ;
            rom[10269] = 8'hf7 ;
            rom[10270] = 8'heb ;
            rom[10271] = 8'h02 ;
            rom[10272] = 8'hec ;
            rom[10273] = 8'hfe ;
            rom[10274] = 8'hd6 ;
            rom[10275] = 8'h0e ;
            rom[10276] = 8'hcc ;
            rom[10277] = 8'hf8 ;
            rom[10278] = 8'h12 ;
            rom[10279] = 8'h0c ;
            rom[10280] = 8'h0b ;
            rom[10281] = 8'hf1 ;
            rom[10282] = 8'h04 ;
            rom[10283] = 8'h26 ;
            rom[10284] = 8'h11 ;
            rom[10285] = 8'hd2 ;
            rom[10286] = 8'hf0 ;
            rom[10287] = 8'h08 ;
            rom[10288] = 8'h11 ;
            rom[10289] = 8'hf9 ;
            rom[10290] = 8'hfd ;
            rom[10291] = 8'h01 ;
            rom[10292] = 8'hed ;
            rom[10293] = 8'h22 ;
            rom[10294] = 8'h19 ;
            rom[10295] = 8'hea ;
            rom[10296] = 8'he3 ;
            rom[10297] = 8'hfd ;
            rom[10298] = 8'h13 ;
            rom[10299] = 8'h02 ;
            rom[10300] = 8'hf3 ;
            rom[10301] = 8'h02 ;
            rom[10302] = 8'h1c ;
            rom[10303] = 8'h13 ;
            rom[10304] = 8'h10 ;
            rom[10305] = 8'h09 ;
            rom[10306] = 8'h23 ;
            rom[10307] = 8'hf9 ;
            rom[10308] = 8'heb ;
            rom[10309] = 8'h02 ;
            rom[10310] = 8'hf5 ;
            rom[10311] = 8'hfc ;
            rom[10312] = 8'hff ;
            rom[10313] = 8'h0c ;
            rom[10314] = 8'he5 ;
            rom[10315] = 8'h04 ;
            rom[10316] = 8'hff ;
            rom[10317] = 8'hee ;
            rom[10318] = 8'h1d ;
            rom[10319] = 8'h17 ;
            rom[10320] = 8'h0c ;
            rom[10321] = 8'hfa ;
            rom[10322] = 8'heb ;
            rom[10323] = 8'hdf ;
            rom[10324] = 8'hd4 ;
            rom[10325] = 8'hdf ;
            rom[10326] = 8'h0d ;
            rom[10327] = 8'h02 ;
            rom[10328] = 8'h31 ;
            rom[10329] = 8'h15 ;
            rom[10330] = 8'h14 ;
            rom[10331] = 8'hf0 ;
            rom[10332] = 8'hef ;
            rom[10333] = 8'hd7 ;
            rom[10334] = 8'h01 ;
            rom[10335] = 8'hee ;
            rom[10336] = 8'h05 ;
            rom[10337] = 8'hf5 ;
            rom[10338] = 8'hee ;
            rom[10339] = 8'hd6 ;
            rom[10340] = 8'hf7 ;
            rom[10341] = 8'hc8 ;
            rom[10342] = 8'h15 ;
            rom[10343] = 8'h19 ;
            rom[10344] = 8'h1d ;
            rom[10345] = 8'h0d ;
            rom[10346] = 8'h14 ;
            rom[10347] = 8'hf8 ;
            rom[10348] = 8'h06 ;
            rom[10349] = 8'hde ;
            rom[10350] = 8'he4 ;
            rom[10351] = 8'hfa ;
            rom[10352] = 8'h25 ;
            rom[10353] = 8'h06 ;
            rom[10354] = 8'h29 ;
            rom[10355] = 8'h00 ;
            rom[10356] = 8'h0c ;
            rom[10357] = 8'h0c ;
            rom[10358] = 8'h04 ;
            rom[10359] = 8'h04 ;
            rom[10360] = 8'h07 ;
            rom[10361] = 8'h0e ;
            rom[10362] = 8'h0e ;
            rom[10363] = 8'he5 ;
            rom[10364] = 8'h13 ;
            rom[10365] = 8'h11 ;
            rom[10366] = 8'hfb ;
            rom[10367] = 8'h0a ;
            rom[10368] = 8'h05 ;
            rom[10369] = 8'he9 ;
            rom[10370] = 8'h16 ;
            rom[10371] = 8'hd8 ;
            rom[10372] = 8'hd7 ;
            rom[10373] = 8'hf3 ;
            rom[10374] = 8'h1b ;
            rom[10375] = 8'h08 ;
            rom[10376] = 8'hc5 ;
            rom[10377] = 8'hf0 ;
            rom[10378] = 8'h0d ;
            rom[10379] = 8'h16 ;
            rom[10380] = 8'hf7 ;
            rom[10381] = 8'he1 ;
            rom[10382] = 8'hf8 ;
            rom[10383] = 8'hfb ;
            rom[10384] = 8'h04 ;
            rom[10385] = 8'h18 ;
            rom[10386] = 8'h19 ;
            rom[10387] = 8'h07 ;
            rom[10388] = 8'he4 ;
            rom[10389] = 8'hff ;
            rom[10390] = 8'h0e ;
            rom[10391] = 8'hda ;
            rom[10392] = 8'hf0 ;
            rom[10393] = 8'h0f ;
            rom[10394] = 8'hfb ;
            rom[10395] = 8'hf6 ;
            rom[10396] = 8'hea ;
            rom[10397] = 8'h03 ;
            rom[10398] = 8'hfa ;
            rom[10399] = 8'h05 ;
            rom[10400] = 8'hf5 ;
            rom[10401] = 8'h02 ;
            rom[10402] = 8'h04 ;
            rom[10403] = 8'hcc ;
            rom[10404] = 8'h03 ;
            rom[10405] = 8'h1d ;
            rom[10406] = 8'hff ;
            rom[10407] = 8'hd7 ;
            rom[10408] = 8'hfa ;
            rom[10409] = 8'hd9 ;
            rom[10410] = 8'h14 ;
            rom[10411] = 8'hf7 ;
            rom[10412] = 8'h18 ;
            rom[10413] = 8'h05 ;
            rom[10414] = 8'hf8 ;
            rom[10415] = 8'he4 ;
            rom[10416] = 8'h03 ;
            rom[10417] = 8'hd4 ;
            rom[10418] = 8'h01 ;
            rom[10419] = 8'h11 ;
            rom[10420] = 8'hcb ;
            rom[10421] = 8'h15 ;
            rom[10422] = 8'h14 ;
            rom[10423] = 8'he5 ;
            rom[10424] = 8'he6 ;
            rom[10425] = 8'hf2 ;
            rom[10426] = 8'h31 ;
            rom[10427] = 8'h00 ;
            rom[10428] = 8'h17 ;
            rom[10429] = 8'h1c ;
            rom[10430] = 8'hf8 ;
            rom[10431] = 8'h02 ;
            rom[10432] = 8'hf8 ;
            rom[10433] = 8'h01 ;
            rom[10434] = 8'h00 ;
            rom[10435] = 8'hea ;
            rom[10436] = 8'hfe ;
            rom[10437] = 8'h35 ;
            rom[10438] = 8'hfe ;
            rom[10439] = 8'h2d ;
            rom[10440] = 8'hf1 ;
            rom[10441] = 8'h08 ;
            rom[10442] = 8'he5 ;
            rom[10443] = 8'h0c ;
            rom[10444] = 8'he0 ;
            rom[10445] = 8'hde ;
            rom[10446] = 8'he6 ;
            rom[10447] = 8'h1d ;
            rom[10448] = 8'he5 ;
            rom[10449] = 8'hf5 ;
            rom[10450] = 8'h1e ;
            rom[10451] = 8'he9 ;
            rom[10452] = 8'hf0 ;
            rom[10453] = 8'hdc ;
            rom[10454] = 8'h13 ;
            rom[10455] = 8'h07 ;
            rom[10456] = 8'h1a ;
            rom[10457] = 8'h11 ;
            rom[10458] = 8'h33 ;
            rom[10459] = 8'hf3 ;
            rom[10460] = 8'hd6 ;
            rom[10461] = 8'hd7 ;
            rom[10462] = 8'h04 ;
            rom[10463] = 8'hfd ;
            rom[10464] = 8'h12 ;
            rom[10465] = 8'h0e ;
            rom[10466] = 8'hea ;
            rom[10467] = 8'h04 ;
            rom[10468] = 8'he8 ;
            rom[10469] = 8'h02 ;
            rom[10470] = 8'h10 ;
            rom[10471] = 8'hfa ;
            rom[10472] = 8'h1c ;
            rom[10473] = 8'h12 ;
            rom[10474] = 8'h0a ;
            rom[10475] = 8'hfd ;
            rom[10476] = 8'hdf ;
            rom[10477] = 8'h0c ;
            rom[10478] = 8'hea ;
            rom[10479] = 8'hfb ;
            rom[10480] = 8'h13 ;
            rom[10481] = 8'hfa ;
            rom[10482] = 8'he4 ;
            rom[10483] = 8'he5 ;
            rom[10484] = 8'he0 ;
            rom[10485] = 8'h2b ;
            rom[10486] = 8'hea ;
            rom[10487] = 8'h08 ;
            rom[10488] = 8'h02 ;
            rom[10489] = 8'hf5 ;
            rom[10490] = 8'h09 ;
            rom[10491] = 8'hff ;
            rom[10492] = 8'h0d ;
            rom[10493] = 8'h0b ;
            rom[10494] = 8'h0c ;
            rom[10495] = 8'hea ;
            rom[10496] = 8'h17 ;
            rom[10497] = 8'hf4 ;
            rom[10498] = 8'h16 ;
            rom[10499] = 8'h14 ;
            rom[10500] = 8'hfd ;
            rom[10501] = 8'h07 ;
            rom[10502] = 8'hdd ;
            rom[10503] = 8'h00 ;
            rom[10504] = 8'h02 ;
            rom[10505] = 8'hf9 ;
            rom[10506] = 8'h1e ;
            rom[10507] = 8'h09 ;
            rom[10508] = 8'h14 ;
            rom[10509] = 8'he9 ;
            rom[10510] = 8'h1c ;
            rom[10511] = 8'h17 ;
            rom[10512] = 8'hec ;
            rom[10513] = 8'hfc ;
            rom[10514] = 8'h04 ;
            rom[10515] = 8'hf7 ;
            rom[10516] = 8'h0a ;
            rom[10517] = 8'heb ;
            rom[10518] = 8'he4 ;
            rom[10519] = 8'hf0 ;
            rom[10520] = 8'he1 ;
            rom[10521] = 8'hf2 ;
            rom[10522] = 8'hf3 ;
            rom[10523] = 8'hf1 ;
            rom[10524] = 8'h04 ;
            rom[10525] = 8'hd6 ;
            rom[10526] = 8'h19 ;
            rom[10527] = 8'hdc ;
            rom[10528] = 8'hce ;
            rom[10529] = 8'h0c ;
            rom[10530] = 8'hf0 ;
            rom[10531] = 8'h0d ;
            rom[10532] = 8'hfd ;
            rom[10533] = 8'h2c ;
            rom[10534] = 8'he9 ;
            rom[10535] = 8'hf6 ;
            rom[10536] = 8'hfe ;
            rom[10537] = 8'hfa ;
            rom[10538] = 8'h06 ;
            rom[10539] = 8'h0f ;
            rom[10540] = 8'hfd ;
            rom[10541] = 8'h18 ;
            rom[10542] = 8'hfc ;
            rom[10543] = 8'hd4 ;
            rom[10544] = 8'he1 ;
            rom[10545] = 8'hd5 ;
            rom[10546] = 8'hec ;
            rom[10547] = 8'h1d ;
            rom[10548] = 8'hf7 ;
            rom[10549] = 8'h11 ;
            rom[10550] = 8'hc9 ;
            rom[10551] = 8'hd4 ;
            rom[10552] = 8'h17 ;
            rom[10553] = 8'hf1 ;
            rom[10554] = 8'h0a ;
            rom[10555] = 8'h33 ;
            rom[10556] = 8'hf3 ;
            rom[10557] = 8'h0d ;
            rom[10558] = 8'h20 ;
            rom[10559] = 8'heb ;
            rom[10560] = 8'hf7 ;
            rom[10561] = 8'h18 ;
            rom[10562] = 8'hf3 ;
            rom[10563] = 8'heb ;
            rom[10564] = 8'hf0 ;
            rom[10565] = 8'h09 ;
            rom[10566] = 8'h02 ;
            rom[10567] = 8'hff ;
            rom[10568] = 8'h32 ;
            rom[10569] = 8'he5 ;
            rom[10570] = 8'hde ;
            rom[10571] = 8'hfa ;
            rom[10572] = 8'hf5 ;
            rom[10573] = 8'hf9 ;
            rom[10574] = 8'h1f ;
            rom[10575] = 8'h18 ;
            rom[10576] = 8'h18 ;
            rom[10577] = 8'h23 ;
            rom[10578] = 8'hfa ;
            rom[10579] = 8'h05 ;
            rom[10580] = 8'h06 ;
            rom[10581] = 8'hcc ;
            rom[10582] = 8'hfe ;
            rom[10583] = 8'he9 ;
            rom[10584] = 8'h1d ;
            rom[10585] = 8'hf6 ;
            rom[10586] = 8'he8 ;
            rom[10587] = 8'h0a ;
            rom[10588] = 8'hf2 ;
            rom[10589] = 8'hea ;
            rom[10590] = 8'h08 ;
            rom[10591] = 8'h25 ;
            rom[10592] = 8'h0b ;
            rom[10593] = 8'h36 ;
            rom[10594] = 8'hd9 ;
            rom[10595] = 8'hf2 ;
            rom[10596] = 8'he5 ;
            rom[10597] = 8'he2 ;
            rom[10598] = 8'h1b ;
            rom[10599] = 8'hff ;
            rom[10600] = 8'hfd ;
            rom[10601] = 8'hfb ;
            rom[10602] = 8'h15 ;
            rom[10603] = 8'he2 ;
            rom[10604] = 8'hfa ;
            rom[10605] = 8'h01 ;
            rom[10606] = 8'h17 ;
            rom[10607] = 8'hff ;
            rom[10608] = 8'hf4 ;
            rom[10609] = 8'he5 ;
            rom[10610] = 8'hfc ;
            rom[10611] = 8'hf4 ;
            rom[10612] = 8'h03 ;
            rom[10613] = 8'h18 ;
            rom[10614] = 8'h0b ;
            rom[10615] = 8'hff ;
            rom[10616] = 8'h0a ;
            rom[10617] = 8'h13 ;
            rom[10618] = 8'h22 ;
            rom[10619] = 8'hea ;
            rom[10620] = 8'hd1 ;
            rom[10621] = 8'he5 ;
            rom[10622] = 8'h1b ;
            rom[10623] = 8'hd2 ;
            rom[10624] = 8'hed ;
            rom[10625] = 8'h10 ;
            rom[10626] = 8'hdb ;
            rom[10627] = 8'hf6 ;
            rom[10628] = 8'hf4 ;
            rom[10629] = 8'h08 ;
            rom[10630] = 8'hff ;
            rom[10631] = 8'h11 ;
            rom[10632] = 8'h20 ;
            rom[10633] = 8'hf5 ;
            rom[10634] = 8'h0f ;
            rom[10635] = 8'h02 ;
            rom[10636] = 8'h04 ;
            rom[10637] = 8'h09 ;
            rom[10638] = 8'h20 ;
            rom[10639] = 8'h18 ;
            rom[10640] = 8'hf7 ;
            rom[10641] = 8'h19 ;
            rom[10642] = 8'h04 ;
            rom[10643] = 8'h0b ;
            rom[10644] = 8'hed ;
            rom[10645] = 8'h0f ;
            rom[10646] = 8'h0b ;
            rom[10647] = 8'h07 ;
            rom[10648] = 8'h0d ;
            rom[10649] = 8'hf1 ;
            rom[10650] = 8'h00 ;
            rom[10651] = 8'he4 ;
            rom[10652] = 8'h03 ;
            rom[10653] = 8'h01 ;
            rom[10654] = 8'hfd ;
            rom[10655] = 8'h16 ;
            rom[10656] = 8'h0d ;
            rom[10657] = 8'hd1 ;
            rom[10658] = 8'hee ;
            rom[10659] = 8'h0a ;
            rom[10660] = 8'hdb ;
            rom[10661] = 8'h0c ;
            rom[10662] = 8'h04 ;
            rom[10663] = 8'h0c ;
            rom[10664] = 8'hff ;
            rom[10665] = 8'h0e ;
            rom[10666] = 8'h03 ;
            rom[10667] = 8'h1d ;
            rom[10668] = 8'h00 ;
            rom[10669] = 8'h07 ;
            rom[10670] = 8'he4 ;
            rom[10671] = 8'h11 ;
            rom[10672] = 8'hdf ;
            rom[10673] = 8'h02 ;
            rom[10674] = 8'hf1 ;
            rom[10675] = 8'h0f ;
            rom[10676] = 8'h19 ;
            rom[10677] = 8'h07 ;
            rom[10678] = 8'h1a ;
            rom[10679] = 8'h13 ;
            rom[10680] = 8'hf5 ;
            rom[10681] = 8'hea ;
            rom[10682] = 8'hfa ;
            rom[10683] = 8'h0c ;
            rom[10684] = 8'h0a ;
            rom[10685] = 8'hf9 ;
            rom[10686] = 8'hfe ;
            rom[10687] = 8'h26 ;
            rom[10688] = 8'h14 ;
            rom[10689] = 8'h08 ;
            rom[10690] = 8'hf4 ;
            rom[10691] = 8'hfb ;
            rom[10692] = 8'h03 ;
            rom[10693] = 8'h12 ;
            rom[10694] = 8'hf5 ;
            rom[10695] = 8'h01 ;
            rom[10696] = 8'h1e ;
            rom[10697] = 8'h28 ;
            rom[10698] = 8'hd1 ;
            rom[10699] = 8'he7 ;
            rom[10700] = 8'h0f ;
            rom[10701] = 8'h0c ;
            rom[10702] = 8'h32 ;
            rom[10703] = 8'he6 ;
            rom[10704] = 8'h1c ;
            rom[10705] = 8'hfe ;
            rom[10706] = 8'h01 ;
            rom[10707] = 8'he1 ;
            rom[10708] = 8'hc1 ;
            rom[10709] = 8'h18 ;
            rom[10710] = 8'hf3 ;
            rom[10711] = 8'hfd ;
            rom[10712] = 8'hea ;
            rom[10713] = 8'h1f ;
            rom[10714] = 8'hf2 ;
            rom[10715] = 8'hfa ;
            rom[10716] = 8'h09 ;
            rom[10717] = 8'hee ;
            rom[10718] = 8'hf7 ;
            rom[10719] = 8'h04 ;
            rom[10720] = 8'h02 ;
            rom[10721] = 8'h19 ;
            rom[10722] = 8'h0e ;
            rom[10723] = 8'hf9 ;
            rom[10724] = 8'hf5 ;
            rom[10725] = 8'hde ;
            rom[10726] = 8'hf7 ;
            rom[10727] = 8'h21 ;
            rom[10728] = 8'h0d ;
            rom[10729] = 8'h23 ;
            rom[10730] = 8'he4 ;
            rom[10731] = 8'h19 ;
            rom[10732] = 8'h1a ;
            rom[10733] = 8'h09 ;
            rom[10734] = 8'hf8 ;
            rom[10735] = 8'h00 ;
            rom[10736] = 8'h00 ;
            rom[10737] = 8'h07 ;
            rom[10738] = 8'h0f ;
            rom[10739] = 8'he7 ;
            rom[10740] = 8'h05 ;
            rom[10741] = 8'he1 ;
            rom[10742] = 8'h0e ;
            rom[10743] = 8'heb ;
            rom[10744] = 8'hd9 ;
            rom[10745] = 8'h1e ;
            rom[10746] = 8'h08 ;
            rom[10747] = 8'h07 ;
            rom[10748] = 8'hff ;
            rom[10749] = 8'h10 ;
            rom[10750] = 8'h11 ;
            rom[10751] = 8'hff ;
            rom[10752] = 8'hf8 ;
            rom[10753] = 8'h07 ;
            rom[10754] = 8'h16 ;
            rom[10755] = 8'h18 ;
            rom[10756] = 8'h19 ;
            rom[10757] = 8'hb1 ;
            rom[10758] = 8'hf1 ;
            rom[10759] = 8'hde ;
            rom[10760] = 8'hf1 ;
            rom[10761] = 8'h16 ;
            rom[10762] = 8'hea ;
            rom[10763] = 8'he3 ;
            rom[10764] = 8'hd6 ;
            rom[10765] = 8'he5 ;
            rom[10766] = 8'hd5 ;
            rom[10767] = 8'hfc ;
            rom[10768] = 8'h02 ;
            rom[10769] = 8'h0f ;
            rom[10770] = 8'hda ;
            rom[10771] = 8'hc5 ;
            rom[10772] = 8'h12 ;
            rom[10773] = 8'hfd ;
            rom[10774] = 8'hd0 ;
            rom[10775] = 8'he0 ;
            rom[10776] = 8'he1 ;
            rom[10777] = 8'h24 ;
            rom[10778] = 8'h02 ;
            rom[10779] = 8'h05 ;
            rom[10780] = 8'hdc ;
            rom[10781] = 8'h14 ;
            rom[10782] = 8'h27 ;
            rom[10783] = 8'h0d ;
            rom[10784] = 8'hef ;
            rom[10785] = 8'h17 ;
            rom[10786] = 8'hf5 ;
            rom[10787] = 8'hf5 ;
            rom[10788] = 8'hee ;
            rom[10789] = 8'hcf ;
            rom[10790] = 8'he5 ;
            rom[10791] = 8'h1b ;
            rom[10792] = 8'h14 ;
            rom[10793] = 8'h06 ;
            rom[10794] = 8'hc4 ;
            rom[10795] = 8'hbe ;
            rom[10796] = 8'h0a ;
            rom[10797] = 8'hd8 ;
            rom[10798] = 8'h08 ;
            rom[10799] = 8'hef ;
            rom[10800] = 8'hf9 ;
            rom[10801] = 8'h0f ;
            rom[10802] = 8'he1 ;
            rom[10803] = 8'he8 ;
            rom[10804] = 8'h12 ;
            rom[10805] = 8'h08 ;
            rom[10806] = 8'hcf ;
            rom[10807] = 8'hfb ;
            rom[10808] = 8'h18 ;
            rom[10809] = 8'h12 ;
            rom[10810] = 8'h11 ;
            rom[10811] = 8'h09 ;
            rom[10812] = 8'hd7 ;
            rom[10813] = 8'hee ;
            rom[10814] = 8'he5 ;
            rom[10815] = 8'hf8 ;
            rom[10816] = 8'hec ;
            rom[10817] = 8'hc7 ;
            rom[10818] = 8'hec ;
            rom[10819] = 8'hfb ;
            rom[10820] = 8'h08 ;
            rom[10821] = 8'h00 ;
            rom[10822] = 8'hef ;
            rom[10823] = 8'hd8 ;
            rom[10824] = 8'hea ;
            rom[10825] = 8'h00 ;
            rom[10826] = 8'h02 ;
            rom[10827] = 8'h12 ;
            rom[10828] = 8'h0d ;
            rom[10829] = 8'hef ;
            rom[10830] = 8'hfd ;
            rom[10831] = 8'h0b ;
            rom[10832] = 8'hf5 ;
            rom[10833] = 8'he1 ;
            rom[10834] = 8'hef ;
            rom[10835] = 8'hf9 ;
            rom[10836] = 8'hec ;
            rom[10837] = 8'h01 ;
            rom[10838] = 8'hfd ;
            rom[10839] = 8'hfc ;
            rom[10840] = 8'h09 ;
            rom[10841] = 8'hf5 ;
            rom[10842] = 8'h02 ;
            rom[10843] = 8'hee ;
            rom[10844] = 8'h13 ;
            rom[10845] = 8'hf6 ;
            rom[10846] = 8'hfb ;
            rom[10847] = 8'hf9 ;
            rom[10848] = 8'hfe ;
            rom[10849] = 8'hb3 ;
            rom[10850] = 8'h14 ;
            rom[10851] = 8'hc4 ;
            rom[10852] = 8'he7 ;
            rom[10853] = 8'hf1 ;
            rom[10854] = 8'hf0 ;
            rom[10855] = 8'hfe ;
            rom[10856] = 8'hd6 ;
            rom[10857] = 8'hee ;
            rom[10858] = 8'hf6 ;
            rom[10859] = 8'hf6 ;
            rom[10860] = 8'hfc ;
            rom[10861] = 8'hdd ;
            rom[10862] = 8'h0c ;
            rom[10863] = 8'hf5 ;
            rom[10864] = 8'hdd ;
            rom[10865] = 8'h0c ;
            rom[10866] = 8'h1a ;
            rom[10867] = 8'hfa ;
            rom[10868] = 8'h09 ;
            rom[10869] = 8'hee ;
            rom[10870] = 8'h07 ;
            rom[10871] = 8'h03 ;
            rom[10872] = 8'hed ;
            rom[10873] = 8'he5 ;
            rom[10874] = 8'hfe ;
            rom[10875] = 8'h07 ;
            rom[10876] = 8'hfc ;
            rom[10877] = 8'he3 ;
            rom[10878] = 8'he2 ;
            rom[10879] = 8'he4 ;
            rom[10880] = 8'he3 ;
            rom[10881] = 8'hf6 ;
            rom[10882] = 8'h06 ;
            rom[10883] = 8'hf2 ;
            rom[10884] = 8'h0f ;
            rom[10885] = 8'hd6 ;
            rom[10886] = 8'h09 ;
            rom[10887] = 8'hf7 ;
            rom[10888] = 8'hff ;
            rom[10889] = 8'hdc ;
            rom[10890] = 8'h04 ;
            rom[10891] = 8'hf2 ;
            rom[10892] = 8'he8 ;
            rom[10893] = 8'h18 ;
            rom[10894] = 8'hfe ;
            rom[10895] = 8'h16 ;
            rom[10896] = 8'h09 ;
            rom[10897] = 8'h01 ;
            rom[10898] = 8'h0b ;
            rom[10899] = 8'hd0 ;
            rom[10900] = 8'hf1 ;
            rom[10901] = 8'he8 ;
            rom[10902] = 8'hfa ;
            rom[10903] = 8'h03 ;
            rom[10904] = 8'h0b ;
            rom[10905] = 8'hfe ;
            rom[10906] = 8'h15 ;
            rom[10907] = 8'h00 ;
            rom[10908] = 8'h0f ;
            rom[10909] = 8'h3f ;
            rom[10910] = 8'he1 ;
            rom[10911] = 8'h19 ;
            rom[10912] = 8'h10 ;
            rom[10913] = 8'he3 ;
            rom[10914] = 8'h0e ;
            rom[10915] = 8'hbc ;
            rom[10916] = 8'h1d ;
            rom[10917] = 8'hf9 ;
            rom[10918] = 8'h17 ;
            rom[10919] = 8'h23 ;
            rom[10920] = 8'h12 ;
            rom[10921] = 8'h00 ;
            rom[10922] = 8'he7 ;
            rom[10923] = 8'h0c ;
            rom[10924] = 8'h15 ;
            rom[10925] = 8'hfe ;
            rom[10926] = 8'he9 ;
            rom[10927] = 8'h01 ;
            rom[10928] = 8'h08 ;
            rom[10929] = 8'h0c ;
            rom[10930] = 8'h12 ;
            rom[10931] = 8'h0d ;
            rom[10932] = 8'hff ;
            rom[10933] = 8'hf8 ;
            rom[10934] = 8'he5 ;
            rom[10935] = 8'he5 ;
            rom[10936] = 8'h15 ;
            rom[10937] = 8'h06 ;
            rom[10938] = 8'h08 ;
            rom[10939] = 8'h11 ;
            rom[10940] = 8'hf2 ;
            rom[10941] = 8'hd3 ;
            rom[10942] = 8'h02 ;
            rom[10943] = 8'h01 ;
            rom[10944] = 8'hfc ;
            rom[10945] = 8'h17 ;
            rom[10946] = 8'h2e ;
            rom[10947] = 8'heb ;
            rom[10948] = 8'he2 ;
            rom[10949] = 8'hf1 ;
            rom[10950] = 8'hef ;
            rom[10951] = 8'h00 ;
            rom[10952] = 8'hb6 ;
            rom[10953] = 8'he6 ;
            rom[10954] = 8'h07 ;
            rom[10955] = 8'h21 ;
            rom[10956] = 8'hf7 ;
            rom[10957] = 8'hc8 ;
            rom[10958] = 8'hf7 ;
            rom[10959] = 8'h08 ;
            rom[10960] = 8'hc5 ;
            rom[10961] = 8'hec ;
            rom[10962] = 8'h15 ;
            rom[10963] = 8'hfe ;
            rom[10964] = 8'h04 ;
            rom[10965] = 8'h05 ;
            rom[10966] = 8'he2 ;
            rom[10967] = 8'hf0 ;
            rom[10968] = 8'h0b ;
            rom[10969] = 8'h1c ;
            rom[10970] = 8'h07 ;
            rom[10971] = 8'h2a ;
            rom[10972] = 8'hf1 ;
            rom[10973] = 8'h13 ;
            rom[10974] = 8'hee ;
            rom[10975] = 8'hf8 ;
            rom[10976] = 8'hf5 ;
            rom[10977] = 8'h16 ;
            rom[10978] = 8'hef ;
            rom[10979] = 8'hec ;
            rom[10980] = 8'h28 ;
            rom[10981] = 8'h0e ;
            rom[10982] = 8'hfd ;
            rom[10983] = 8'hec ;
            rom[10984] = 8'hfe ;
            rom[10985] = 8'hf7 ;
            rom[10986] = 8'h17 ;
            rom[10987] = 8'h19 ;
            rom[10988] = 8'hac ;
            rom[10989] = 8'h20 ;
            rom[10990] = 8'hde ;
            rom[10991] = 8'h16 ;
            rom[10992] = 8'hf6 ;
            rom[10993] = 8'h1a ;
            rom[10994] = 8'hfa ;
            rom[10995] = 8'h2f ;
            rom[10996] = 8'h13 ;
            rom[10997] = 8'hee ;
            rom[10998] = 8'hf5 ;
            rom[10999] = 8'hf0 ;
            rom[11000] = 8'h1f ;
            rom[11001] = 8'hfe ;
            rom[11002] = 8'h1d ;
            rom[11003] = 8'hf4 ;
            rom[11004] = 8'hf9 ;
            rom[11005] = 8'hf8 ;
            rom[11006] = 8'h09 ;
            rom[11007] = 8'h20 ;
            rom[11008] = 8'h13 ;
            rom[11009] = 8'hff ;
            rom[11010] = 8'hf5 ;
            rom[11011] = 8'h24 ;
            rom[11012] = 8'hff ;
            rom[11013] = 8'hc3 ;
            rom[11014] = 8'h00 ;
            rom[11015] = 8'he7 ;
            rom[11016] = 8'h08 ;
            rom[11017] = 8'hf6 ;
            rom[11018] = 8'he1 ;
            rom[11019] = 8'hfe ;
            rom[11020] = 8'h02 ;
            rom[11021] = 8'h14 ;
            rom[11022] = 8'hcf ;
            rom[11023] = 8'h08 ;
            rom[11024] = 8'hfc ;
            rom[11025] = 8'hf5 ;
            rom[11026] = 8'hf6 ;
            rom[11027] = 8'he2 ;
            rom[11028] = 8'h02 ;
            rom[11029] = 8'h1b ;
            rom[11030] = 8'hfd ;
            rom[11031] = 8'hf3 ;
            rom[11032] = 8'hee ;
            rom[11033] = 8'hf8 ;
            rom[11034] = 8'he8 ;
            rom[11035] = 8'h0e ;
            rom[11036] = 8'hf7 ;
            rom[11037] = 8'hfb ;
            rom[11038] = 8'h06 ;
            rom[11039] = 8'hd1 ;
            rom[11040] = 8'hff ;
            rom[11041] = 8'hf7 ;
            rom[11042] = 8'hd1 ;
            rom[11043] = 8'h0e ;
            rom[11044] = 8'hf8 ;
            rom[11045] = 8'he6 ;
            rom[11046] = 8'h18 ;
            rom[11047] = 8'hfc ;
            rom[11048] = 8'hb9 ;
            rom[11049] = 8'hf1 ;
            rom[11050] = 8'h01 ;
            rom[11051] = 8'h11 ;
            rom[11052] = 8'hea ;
            rom[11053] = 8'hda ;
            rom[11054] = 8'he4 ;
            rom[11055] = 8'h0c ;
            rom[11056] = 8'h06 ;
            rom[11057] = 8'h12 ;
            rom[11058] = 8'he5 ;
            rom[11059] = 8'hf9 ;
            rom[11060] = 8'h10 ;
            rom[11061] = 8'hfd ;
            rom[11062] = 8'hdb ;
            rom[11063] = 8'hf5 ;
            rom[11064] = 8'h21 ;
            rom[11065] = 8'h14 ;
            rom[11066] = 8'heb ;
            rom[11067] = 8'hf3 ;
            rom[11068] = 8'he8 ;
            rom[11069] = 8'h0f ;
            rom[11070] = 8'he6 ;
            rom[11071] = 8'hcd ;
            rom[11072] = 8'h0a ;
            rom[11073] = 8'hea ;
            rom[11074] = 8'he4 ;
            rom[11075] = 8'hf3 ;
            rom[11076] = 8'h0b ;
            rom[11077] = 8'he7 ;
            rom[11078] = 8'he5 ;
            rom[11079] = 8'he4 ;
            rom[11080] = 8'he3 ;
            rom[11081] = 8'he9 ;
            rom[11082] = 8'h09 ;
            rom[11083] = 8'hde ;
            rom[11084] = 8'hfe ;
            rom[11085] = 8'h06 ;
            rom[11086] = 8'hf7 ;
            rom[11087] = 8'hfb ;
            rom[11088] = 8'h04 ;
            rom[11089] = 8'h08 ;
            rom[11090] = 8'hea ;
            rom[11091] = 8'h08 ;
            rom[11092] = 8'h0b ;
            rom[11093] = 8'hd1 ;
            rom[11094] = 8'he4 ;
            rom[11095] = 8'h11 ;
            rom[11096] = 8'h17 ;
            rom[11097] = 8'hf3 ;
            rom[11098] = 8'he7 ;
            rom[11099] = 8'h04 ;
            rom[11100] = 8'he7 ;
            rom[11101] = 8'h08 ;
            rom[11102] = 8'hef ;
            rom[11103] = 8'hdf ;
            rom[11104] = 8'h09 ;
            rom[11105] = 8'he8 ;
            rom[11106] = 8'hd1 ;
            rom[11107] = 8'h07 ;
            rom[11108] = 8'h0a ;
            rom[11109] = 8'h0d ;
            rom[11110] = 8'hf2 ;
            rom[11111] = 8'h01 ;
            rom[11112] = 8'hce ;
            rom[11113] = 8'he9 ;
            rom[11114] = 8'hdd ;
            rom[11115] = 8'hf7 ;
            rom[11116] = 8'hf2 ;
            rom[11117] = 8'h1b ;
            rom[11118] = 8'hef ;
            rom[11119] = 8'h03 ;
            rom[11120] = 8'hfa ;
            rom[11121] = 8'hfe ;
            rom[11122] = 8'hfc ;
            rom[11123] = 8'h18 ;
            rom[11124] = 8'hf9 ;
            rom[11125] = 8'h0a ;
            rom[11126] = 8'hc7 ;
            rom[11127] = 8'hdd ;
            rom[11128] = 8'h15 ;
            rom[11129] = 8'h0c ;
            rom[11130] = 8'hc7 ;
            rom[11131] = 8'h0a ;
            rom[11132] = 8'h01 ;
            rom[11133] = 8'he3 ;
            rom[11134] = 8'hfb ;
            rom[11135] = 8'hfe ;
            rom[11136] = 8'hd9 ;
            rom[11137] = 8'h15 ;
            rom[11138] = 8'he2 ;
            rom[11139] = 8'h02 ;
            rom[11140] = 8'hc4 ;
            rom[11141] = 8'he5 ;
            rom[11142] = 8'h0e ;
            rom[11143] = 8'h1c ;
            rom[11144] = 8'he5 ;
            rom[11145] = 8'hf6 ;
            rom[11146] = 8'he1 ;
            rom[11147] = 8'hf0 ;
            rom[11148] = 8'hf5 ;
            rom[11149] = 8'h06 ;
            rom[11150] = 8'h0d ;
            rom[11151] = 8'hfb ;
            rom[11152] = 8'h00 ;
            rom[11153] = 8'hed ;
            rom[11154] = 8'hd4 ;
            rom[11155] = 8'hfb ;
            rom[11156] = 8'h17 ;
            rom[11157] = 8'hfe ;
            rom[11158] = 8'he2 ;
            rom[11159] = 8'hfe ;
            rom[11160] = 8'hff ;
            rom[11161] = 8'h35 ;
            rom[11162] = 8'hfa ;
            rom[11163] = 8'he6 ;
            rom[11164] = 8'hf6 ;
            rom[11165] = 8'h22 ;
            rom[11166] = 8'hfa ;
            rom[11167] = 8'h0b ;
            rom[11168] = 8'hfe ;
            rom[11169] = 8'hbe ;
            rom[11170] = 8'h26 ;
            rom[11171] = 8'h00 ;
            rom[11172] = 8'h04 ;
            rom[11173] = 8'heb ;
            rom[11174] = 8'h06 ;
            rom[11175] = 8'hda ;
            rom[11176] = 8'hd5 ;
            rom[11177] = 8'hdc ;
            rom[11178] = 8'h1d ;
            rom[11179] = 8'he4 ;
            rom[11180] = 8'h19 ;
            rom[11181] = 8'he1 ;
            rom[11182] = 8'hd7 ;
            rom[11183] = 8'h0f ;
            rom[11184] = 8'h21 ;
            rom[11185] = 8'hf0 ;
            rom[11186] = 8'h19 ;
            rom[11187] = 8'hf7 ;
            rom[11188] = 8'hf0 ;
            rom[11189] = 8'h01 ;
            rom[11190] = 8'hef ;
            rom[11191] = 8'he1 ;
            rom[11192] = 8'hec ;
            rom[11193] = 8'h1f ;
            rom[11194] = 8'h08 ;
            rom[11195] = 8'hf0 ;
            rom[11196] = 8'h07 ;
            rom[11197] = 8'hcb ;
            rom[11198] = 8'h08 ;
            rom[11199] = 8'h18 ;
            rom[11200] = 8'hfd ;
            rom[11201] = 8'h21 ;
            rom[11202] = 8'h08 ;
            rom[11203] = 8'hed ;
            rom[11204] = 8'h05 ;
            rom[11205] = 8'h0e ;
            rom[11206] = 8'h04 ;
            rom[11207] = 8'h05 ;
            rom[11208] = 8'hcb ;
            rom[11209] = 8'h1a ;
            rom[11210] = 8'hd0 ;
            rom[11211] = 8'h01 ;
            rom[11212] = 8'h0e ;
            rom[11213] = 8'hdc ;
            rom[11214] = 8'h06 ;
            rom[11215] = 8'h27 ;
            rom[11216] = 8'hf0 ;
            rom[11217] = 8'h08 ;
            rom[11218] = 8'hf2 ;
            rom[11219] = 8'hf4 ;
            rom[11220] = 8'hd9 ;
            rom[11221] = 8'h0d ;
            rom[11222] = 8'h02 ;
            rom[11223] = 8'hf4 ;
            rom[11224] = 8'h07 ;
            rom[11225] = 8'hf3 ;
            rom[11226] = 8'h32 ;
            rom[11227] = 8'hee ;
            rom[11228] = 8'h06 ;
            rom[11229] = 8'h12 ;
            rom[11230] = 8'hef ;
            rom[11231] = 8'hf8 ;
            rom[11232] = 8'hed ;
            rom[11233] = 8'h28 ;
            rom[11234] = 8'h0c ;
            rom[11235] = 8'h07 ;
            rom[11236] = 8'hed ;
            rom[11237] = 8'h34 ;
            rom[11238] = 8'h10 ;
            rom[11239] = 8'h06 ;
            rom[11240] = 8'h05 ;
            rom[11241] = 8'hfe ;
            rom[11242] = 8'h2a ;
            rom[11243] = 8'h09 ;
            rom[11244] = 8'h14 ;
            rom[11245] = 8'h13 ;
            rom[11246] = 8'hc1 ;
            rom[11247] = 8'he4 ;
            rom[11248] = 8'h19 ;
            rom[11249] = 8'hf4 ;
            rom[11250] = 8'hf6 ;
            rom[11251] = 8'hde ;
            rom[11252] = 8'h17 ;
            rom[11253] = 8'h23 ;
            rom[11254] = 8'h06 ;
            rom[11255] = 8'hf8 ;
            rom[11256] = 8'hf2 ;
            rom[11257] = 8'hf8 ;
            rom[11258] = 8'he8 ;
            rom[11259] = 8'hd2 ;
            rom[11260] = 8'h08 ;
            rom[11261] = 8'h0f ;
            rom[11262] = 8'hff ;
            rom[11263] = 8'h17 ;
            rom[11264] = 8'hd5 ;
            rom[11265] = 8'he7 ;
            rom[11266] = 8'hff ;
            rom[11267] = 8'he8 ;
            rom[11268] = 8'h19 ;
            rom[11269] = 8'h09 ;
            rom[11270] = 8'h03 ;
            rom[11271] = 8'hfa ;
            rom[11272] = 8'h03 ;
            rom[11273] = 8'he0 ;
            rom[11274] = 8'h16 ;
            rom[11275] = 8'h0f ;
            rom[11276] = 8'hff ;
            rom[11277] = 8'hd5 ;
            rom[11278] = 8'h03 ;
            rom[11279] = 8'h2c ;
            rom[11280] = 8'h11 ;
            rom[11281] = 8'hec ;
            rom[11282] = 8'hf5 ;
            rom[11283] = 8'h05 ;
            rom[11284] = 8'hf9 ;
            rom[11285] = 8'hee ;
            rom[11286] = 8'he6 ;
            rom[11287] = 8'hf4 ;
            rom[11288] = 8'h11 ;
            rom[11289] = 8'he9 ;
            rom[11290] = 8'hf9 ;
            rom[11291] = 8'h20 ;
            rom[11292] = 8'hfc ;
            rom[11293] = 8'h1b ;
            rom[11294] = 8'hd6 ;
            rom[11295] = 8'h1b ;
            rom[11296] = 8'hfa ;
            rom[11297] = 8'he7 ;
            rom[11298] = 8'h22 ;
            rom[11299] = 8'h17 ;
            rom[11300] = 8'h16 ;
            rom[11301] = 8'h19 ;
            rom[11302] = 8'h14 ;
            rom[11303] = 8'h07 ;
            rom[11304] = 8'h0e ;
            rom[11305] = 8'h03 ;
            rom[11306] = 8'hfd ;
            rom[11307] = 8'h12 ;
            rom[11308] = 8'h1c ;
            rom[11309] = 8'h1c ;
            rom[11310] = 8'h11 ;
            rom[11311] = 8'hd3 ;
            rom[11312] = 8'h04 ;
            rom[11313] = 8'h03 ;
            rom[11314] = 8'hed ;
            rom[11315] = 8'h15 ;
            rom[11316] = 8'h04 ;
            rom[11317] = 8'h05 ;
            rom[11318] = 8'h04 ;
            rom[11319] = 8'h07 ;
            rom[11320] = 8'h04 ;
            rom[11321] = 8'heb ;
            rom[11322] = 8'h1b ;
            rom[11323] = 8'h09 ;
            rom[11324] = 8'h11 ;
            rom[11325] = 8'h0a ;
            rom[11326] = 8'h01 ;
            rom[11327] = 8'hfb ;
            rom[11328] = 8'hf6 ;
            rom[11329] = 8'h17 ;
            rom[11330] = 8'hf1 ;
            rom[11331] = 8'hfc ;
            rom[11332] = 8'heb ;
            rom[11333] = 8'h00 ;
            rom[11334] = 8'h1b ;
            rom[11335] = 8'h0b ;
            rom[11336] = 8'hff ;
            rom[11337] = 8'h05 ;
            rom[11338] = 8'hda ;
            rom[11339] = 8'hce ;
            rom[11340] = 8'hf6 ;
            rom[11341] = 8'hf3 ;
            rom[11342] = 8'h17 ;
            rom[11343] = 8'hfa ;
            rom[11344] = 8'h0d ;
            rom[11345] = 8'h13 ;
            rom[11346] = 8'he9 ;
            rom[11347] = 8'he1 ;
            rom[11348] = 8'hfd ;
            rom[11349] = 8'h07 ;
            rom[11350] = 8'hf8 ;
            rom[11351] = 8'hcb ;
            rom[11352] = 8'h20 ;
            rom[11353] = 8'hf9 ;
            rom[11354] = 8'h00 ;
            rom[11355] = 8'h1a ;
            rom[11356] = 8'hf0 ;
            rom[11357] = 8'h0e ;
            rom[11358] = 8'hfb ;
            rom[11359] = 8'h25 ;
            rom[11360] = 8'h04 ;
            rom[11361] = 8'h1d ;
            rom[11362] = 8'hf5 ;
            rom[11363] = 8'he2 ;
            rom[11364] = 8'h00 ;
            rom[11365] = 8'h09 ;
            rom[11366] = 8'h01 ;
            rom[11367] = 8'h10 ;
            rom[11368] = 8'h10 ;
            rom[11369] = 8'h02 ;
            rom[11370] = 8'h24 ;
            rom[11371] = 8'h0d ;
            rom[11372] = 8'hf8 ;
            rom[11373] = 8'hcb ;
            rom[11374] = 8'hee ;
            rom[11375] = 8'hf9 ;
            rom[11376] = 8'hcd ;
            rom[11377] = 8'hfb ;
            rom[11378] = 8'h1f ;
            rom[11379] = 8'h11 ;
            rom[11380] = 8'h2d ;
            rom[11381] = 8'h0d ;
            rom[11382] = 8'h16 ;
            rom[11383] = 8'hfa ;
            rom[11384] = 8'h07 ;
            rom[11385] = 8'h04 ;
            rom[11386] = 8'h09 ;
            rom[11387] = 8'hff ;
            rom[11388] = 8'he4 ;
            rom[11389] = 8'hfa ;
            rom[11390] = 8'h14 ;
            rom[11391] = 8'he0 ;
            rom[11392] = 8'hca ;
            rom[11393] = 8'h24 ;
            rom[11394] = 8'h03 ;
            rom[11395] = 8'hfd ;
            rom[11396] = 8'hcb ;
            rom[11397] = 8'h09 ;
            rom[11398] = 8'h0a ;
            rom[11399] = 8'hd5 ;
            rom[11400] = 8'hf9 ;
            rom[11401] = 8'h01 ;
            rom[11402] = 8'h16 ;
            rom[11403] = 8'hf7 ;
            rom[11404] = 8'he8 ;
            rom[11405] = 8'h00 ;
            rom[11406] = 8'hf9 ;
            rom[11407] = 8'h11 ;
            rom[11408] = 8'hf8 ;
            rom[11409] = 8'he2 ;
            rom[11410] = 8'h22 ;
            rom[11411] = 8'hd3 ;
            rom[11412] = 8'hfc ;
            rom[11413] = 8'h03 ;
            rom[11414] = 8'h01 ;
            rom[11415] = 8'hf4 ;
            rom[11416] = 8'hfd ;
            rom[11417] = 8'h2d ;
            rom[11418] = 8'hee ;
            rom[11419] = 8'h03 ;
            rom[11420] = 8'h07 ;
            rom[11421] = 8'hf1 ;
            rom[11422] = 8'h02 ;
            rom[11423] = 8'hbd ;
            rom[11424] = 8'hd5 ;
            rom[11425] = 8'hdd ;
            rom[11426] = 8'h12 ;
            rom[11427] = 8'hde ;
            rom[11428] = 8'ha7 ;
            rom[11429] = 8'h03 ;
            rom[11430] = 8'hfa ;
            rom[11431] = 8'h02 ;
            rom[11432] = 8'hf5 ;
            rom[11433] = 8'hd9 ;
            rom[11434] = 8'hf6 ;
            rom[11435] = 8'h18 ;
            rom[11436] = 8'h2f ;
            rom[11437] = 8'he3 ;
            rom[11438] = 8'h08 ;
            rom[11439] = 8'hff ;
            rom[11440] = 8'he6 ;
            rom[11441] = 8'hf4 ;
            rom[11442] = 8'h00 ;
            rom[11443] = 8'h18 ;
            rom[11444] = 8'h0a ;
            rom[11445] = 8'hf8 ;
            rom[11446] = 8'h00 ;
            rom[11447] = 8'h13 ;
            rom[11448] = 8'hfe ;
            rom[11449] = 8'he9 ;
            rom[11450] = 8'h04 ;
            rom[11451] = 8'he8 ;
            rom[11452] = 8'h09 ;
            rom[11453] = 8'he4 ;
            rom[11454] = 8'h11 ;
            rom[11455] = 8'h14 ;
            rom[11456] = 8'h17 ;
            rom[11457] = 8'he7 ;
            rom[11458] = 8'h11 ;
            rom[11459] = 8'h0a ;
            rom[11460] = 8'he2 ;
            rom[11461] = 8'h0f ;
            rom[11462] = 8'h18 ;
            rom[11463] = 8'hfd ;
            rom[11464] = 8'hfe ;
            rom[11465] = 8'hf2 ;
            rom[11466] = 8'hfb ;
            rom[11467] = 8'hf3 ;
            rom[11468] = 8'h07 ;
            rom[11469] = 8'hdc ;
            rom[11470] = 8'hec ;
            rom[11471] = 8'h03 ;
            rom[11472] = 8'h03 ;
            rom[11473] = 8'hf2 ;
            rom[11474] = 8'hf7 ;
            rom[11475] = 8'hd5 ;
            rom[11476] = 8'hde ;
            rom[11477] = 8'hed ;
            rom[11478] = 8'hde ;
            rom[11479] = 8'h0b ;
            rom[11480] = 8'h06 ;
            rom[11481] = 8'h0f ;
            rom[11482] = 8'he7 ;
            rom[11483] = 8'hec ;
            rom[11484] = 8'he4 ;
            rom[11485] = 8'hfc ;
            rom[11486] = 8'hd7 ;
            rom[11487] = 8'h0b ;
            rom[11488] = 8'hff ;
            rom[11489] = 8'h19 ;
            rom[11490] = 8'he4 ;
            rom[11491] = 8'h06 ;
            rom[11492] = 8'h00 ;
            rom[11493] = 8'hee ;
            rom[11494] = 8'hed ;
            rom[11495] = 8'h01 ;
            rom[11496] = 8'h00 ;
            rom[11497] = 8'he0 ;
            rom[11498] = 8'h09 ;
            rom[11499] = 8'he6 ;
            rom[11500] = 8'h0e ;
            rom[11501] = 8'h02 ;
            rom[11502] = 8'h04 ;
            rom[11503] = 8'h05 ;
            rom[11504] = 8'h21 ;
            rom[11505] = 8'hdc ;
            rom[11506] = 8'h14 ;
            rom[11507] = 8'h14 ;
            rom[11508] = 8'h2e ;
            rom[11509] = 8'hf3 ;
            rom[11510] = 8'h02 ;
            rom[11511] = 8'hf3 ;
            rom[11512] = 8'hf9 ;
            rom[11513] = 8'hf0 ;
            rom[11514] = 8'h08 ;
            rom[11515] = 8'hee ;
            rom[11516] = 8'hfb ;
            rom[11517] = 8'hf2 ;
            rom[11518] = 8'hfc ;
            rom[11519] = 8'hf3 ;
            rom[11520] = 8'hd9 ;
            rom[11521] = 8'hf1 ;
            rom[11522] = 8'h0f ;
            rom[11523] = 8'hfd ;
            rom[11524] = 8'h01 ;
            rom[11525] = 8'hf1 ;
            rom[11526] = 8'hd8 ;
            rom[11527] = 8'h09 ;
            rom[11528] = 8'hff ;
            rom[11529] = 8'h01 ;
            rom[11530] = 8'hf1 ;
            rom[11531] = 8'hff ;
            rom[11532] = 8'hd5 ;
            rom[11533] = 8'hdf ;
            rom[11534] = 8'h18 ;
            rom[11535] = 8'h17 ;
            rom[11536] = 8'h07 ;
            rom[11537] = 8'h07 ;
            rom[11538] = 8'h1f ;
            rom[11539] = 8'h2a ;
            rom[11540] = 8'hf0 ;
            rom[11541] = 8'hfb ;
            rom[11542] = 8'h03 ;
            rom[11543] = 8'h28 ;
            rom[11544] = 8'h26 ;
            rom[11545] = 8'hbf ;
            rom[11546] = 8'hf5 ;
            rom[11547] = 8'hd7 ;
            rom[11548] = 8'hff ;
            rom[11549] = 8'h1b ;
            rom[11550] = 8'h15 ;
            rom[11551] = 8'h18 ;
            rom[11552] = 8'h04 ;
            rom[11553] = 8'h00 ;
            rom[11554] = 8'h17 ;
            rom[11555] = 8'hec ;
            rom[11556] = 8'h2e ;
            rom[11557] = 8'hf0 ;
            rom[11558] = 8'hf3 ;
            rom[11559] = 8'he7 ;
            rom[11560] = 8'he6 ;
            rom[11561] = 8'h00 ;
            rom[11562] = 8'he3 ;
            rom[11563] = 8'h17 ;
            rom[11564] = 8'h02 ;
            rom[11565] = 8'h11 ;
            rom[11566] = 8'h02 ;
            rom[11567] = 8'hf0 ;
            rom[11568] = 8'h06 ;
            rom[11569] = 8'hd8 ;
            rom[11570] = 8'h06 ;
            rom[11571] = 8'hf0 ;
            rom[11572] = 8'hec ;
            rom[11573] = 8'h0d ;
            rom[11574] = 8'he3 ;
            rom[11575] = 8'h0d ;
            rom[11576] = 8'h03 ;
            rom[11577] = 8'h0e ;
            rom[11578] = 8'hfe ;
            rom[11579] = 8'hdf ;
            rom[11580] = 8'h10 ;
            rom[11581] = 8'hd4 ;
            rom[11582] = 8'h23 ;
            rom[11583] = 8'h06 ;
            rom[11584] = 8'hed ;
            rom[11585] = 8'h37 ;
            rom[11586] = 8'h1b ;
            rom[11587] = 8'h15 ;
            rom[11588] = 8'h02 ;
            rom[11589] = 8'h12 ;
            rom[11590] = 8'hdf ;
            rom[11591] = 8'h03 ;
            rom[11592] = 8'hcd ;
            rom[11593] = 8'h13 ;
            rom[11594] = 8'hf4 ;
            rom[11595] = 8'hf8 ;
            rom[11596] = 8'hfa ;
            rom[11597] = 8'h15 ;
            rom[11598] = 8'he5 ;
            rom[11599] = 8'h20 ;
            rom[11600] = 8'hff ;
            rom[11601] = 8'h01 ;
            rom[11602] = 8'hf2 ;
            rom[11603] = 8'hed ;
            rom[11604] = 8'h0c ;
            rom[11605] = 8'h13 ;
            rom[11606] = 8'h05 ;
            rom[11607] = 8'hec ;
            rom[11608] = 8'hda ;
            rom[11609] = 8'h1f ;
            rom[11610] = 8'h04 ;
            rom[11611] = 8'hfe ;
            rom[11612] = 8'heb ;
            rom[11613] = 8'h06 ;
            rom[11614] = 8'hee ;
            rom[11615] = 8'h03 ;
            rom[11616] = 8'h1a ;
            rom[11617] = 8'hf9 ;
            rom[11618] = 8'hfa ;
            rom[11619] = 8'h00 ;
            rom[11620] = 8'hf0 ;
            rom[11621] = 8'h08 ;
            rom[11622] = 8'h05 ;
            rom[11623] = 8'hfa ;
            rom[11624] = 8'hff ;
            rom[11625] = 8'hf1 ;
            rom[11626] = 8'he9 ;
            rom[11627] = 8'h32 ;
            rom[11628] = 8'hf1 ;
            rom[11629] = 8'hdf ;
            rom[11630] = 8'h10 ;
            rom[11631] = 8'hf3 ;
            rom[11632] = 8'h06 ;
            rom[11633] = 8'h0d ;
            rom[11634] = 8'hf2 ;
            rom[11635] = 8'h06 ;
            rom[11636] = 8'h38 ;
            rom[11637] = 8'h12 ;
            rom[11638] = 8'h01 ;
            rom[11639] = 8'hd7 ;
            rom[11640] = 8'h00 ;
            rom[11641] = 8'h38 ;
            rom[11642] = 8'h0c ;
            rom[11643] = 8'h02 ;
            rom[11644] = 8'hfd ;
            rom[11645] = 8'h00 ;
            rom[11646] = 8'hfd ;
            rom[11647] = 8'h1c ;
            rom[11648] = 8'hdd ;
            rom[11649] = 8'h17 ;
            rom[11650] = 8'hf0 ;
            rom[11651] = 8'hfc ;
            rom[11652] = 8'h0a ;
            rom[11653] = 8'hd4 ;
            rom[11654] = 8'he8 ;
            rom[11655] = 8'he8 ;
            rom[11656] = 8'hfa ;
            rom[11657] = 8'hec ;
            rom[11658] = 8'h15 ;
            rom[11659] = 8'hc3 ;
            rom[11660] = 8'he9 ;
            rom[11661] = 8'h07 ;
            rom[11662] = 8'hfe ;
            rom[11663] = 8'hb5 ;
            rom[11664] = 8'he8 ;
            rom[11665] = 8'h03 ;
            rom[11666] = 8'h09 ;
            rom[11667] = 8'hfa ;
            rom[11668] = 8'hda ;
            rom[11669] = 8'hff ;
            rom[11670] = 8'h19 ;
            rom[11671] = 8'hdb ;
            rom[11672] = 8'h02 ;
            rom[11673] = 8'h05 ;
            rom[11674] = 8'h03 ;
            rom[11675] = 8'h0d ;
            rom[11676] = 8'h0b ;
            rom[11677] = 8'hff ;
            rom[11678] = 8'h0d ;
            rom[11679] = 8'h23 ;
            rom[11680] = 8'h08 ;
            rom[11681] = 8'h03 ;
            rom[11682] = 8'hf0 ;
            rom[11683] = 8'h0f ;
            rom[11684] = 8'h08 ;
            rom[11685] = 8'hea ;
            rom[11686] = 8'hed ;
            rom[11687] = 8'h24 ;
            rom[11688] = 8'hea ;
            rom[11689] = 8'he4 ;
            rom[11690] = 8'he6 ;
            rom[11691] = 8'hf9 ;
            rom[11692] = 8'heb ;
            rom[11693] = 8'he3 ;
            rom[11694] = 8'hf1 ;
            rom[11695] = 8'h0d ;
            rom[11696] = 8'h0a ;
            rom[11697] = 8'h22 ;
            rom[11698] = 8'hf3 ;
            rom[11699] = 8'hf8 ;
            rom[11700] = 8'hf7 ;
            rom[11701] = 8'h18 ;
            rom[11702] = 8'h07 ;
            rom[11703] = 8'h03 ;
            rom[11704] = 8'h18 ;
            rom[11705] = 8'hed ;
            rom[11706] = 8'h04 ;
            rom[11707] = 8'h0e ;
            rom[11708] = 8'h24 ;
            rom[11709] = 8'he0 ;
            rom[11710] = 8'hea ;
            rom[11711] = 8'hf2 ;
            rom[11712] = 8'h1b ;
            rom[11713] = 8'h00 ;
            rom[11714] = 8'h21 ;
            rom[11715] = 8'he8 ;
            rom[11716] = 8'h0c ;
            rom[11717] = 8'h29 ;
            rom[11718] = 8'hdf ;
            rom[11719] = 8'h00 ;
            rom[11720] = 8'hf7 ;
            rom[11721] = 8'hfa ;
            rom[11722] = 8'hcf ;
            rom[11723] = 8'he6 ;
            rom[11724] = 8'hdf ;
            rom[11725] = 8'he8 ;
            rom[11726] = 8'he7 ;
            rom[11727] = 8'h12 ;
            rom[11728] = 8'h23 ;
            rom[11729] = 8'hef ;
            rom[11730] = 8'hea ;
            rom[11731] = 8'hfb ;
            rom[11732] = 8'hfc ;
            rom[11733] = 8'he4 ;
            rom[11734] = 8'he1 ;
            rom[11735] = 8'h05 ;
            rom[11736] = 8'hfd ;
            rom[11737] = 8'h13 ;
            rom[11738] = 8'he6 ;
            rom[11739] = 8'hef ;
            rom[11740] = 8'hb7 ;
            rom[11741] = 8'hf8 ;
            rom[11742] = 8'hc3 ;
            rom[11743] = 8'hb3 ;
            rom[11744] = 8'he9 ;
            rom[11745] = 8'h00 ;
            rom[11746] = 8'h03 ;
            rom[11747] = 8'hfd ;
            rom[11748] = 8'hf5 ;
            rom[11749] = 8'h0f ;
            rom[11750] = 8'h1d ;
            rom[11751] = 8'h01 ;
            rom[11752] = 8'he9 ;
            rom[11753] = 8'h12 ;
            rom[11754] = 8'h13 ;
            rom[11755] = 8'hed ;
            rom[11756] = 8'hf9 ;
            rom[11757] = 8'h15 ;
            rom[11758] = 8'hf3 ;
            rom[11759] = 8'h08 ;
            rom[11760] = 8'hf8 ;
            rom[11761] = 8'hea ;
            rom[11762] = 8'h19 ;
            rom[11763] = 8'hd1 ;
            rom[11764] = 8'h00 ;
            rom[11765] = 8'hec ;
            rom[11766] = 8'h0c ;
            rom[11767] = 8'h27 ;
            rom[11768] = 8'he1 ;
            rom[11769] = 8'hf9 ;
            rom[11770] = 8'hcf ;
            rom[11771] = 8'h03 ;
            rom[11772] = 8'hd2 ;
            rom[11773] = 8'h12 ;
            rom[11774] = 8'h03 ;
            rom[11775] = 8'hec ;
            rom[11776] = 8'h0a ;
            rom[11777] = 8'hdf ;
            rom[11778] = 8'h17 ;
            rom[11779] = 8'hca ;
            rom[11780] = 8'he5 ;
            rom[11781] = 8'h1c ;
            rom[11782] = 8'hfe ;
            rom[11783] = 8'hd4 ;
            rom[11784] = 8'h00 ;
            rom[11785] = 8'h00 ;
            rom[11786] = 8'h01 ;
            rom[11787] = 8'h17 ;
            rom[11788] = 8'hee ;
            rom[11789] = 8'hff ;
            rom[11790] = 8'h19 ;
            rom[11791] = 8'hf7 ;
            rom[11792] = 8'hf4 ;
            rom[11793] = 8'h1a ;
            rom[11794] = 8'hff ;
            rom[11795] = 8'hf9 ;
            rom[11796] = 8'he2 ;
            rom[11797] = 8'hc5 ;
            rom[11798] = 8'h14 ;
            rom[11799] = 8'h0b ;
            rom[11800] = 8'hd3 ;
            rom[11801] = 8'he1 ;
            rom[11802] = 8'hf4 ;
            rom[11803] = 8'hb4 ;
            rom[11804] = 8'he0 ;
            rom[11805] = 8'hdd ;
            rom[11806] = 8'hd1 ;
            rom[11807] = 8'hff ;
            rom[11808] = 8'he5 ;
            rom[11809] = 8'h0a ;
            rom[11810] = 8'h1a ;
            rom[11811] = 8'h03 ;
            rom[11812] = 8'h10 ;
            rom[11813] = 8'he7 ;
            rom[11814] = 8'h05 ;
            rom[11815] = 8'hc7 ;
            rom[11816] = 8'h16 ;
            rom[11817] = 8'hf8 ;
            rom[11818] = 8'hff ;
            rom[11819] = 8'h11 ;
            rom[11820] = 8'h00 ;
            rom[11821] = 8'he6 ;
            rom[11822] = 8'h01 ;
            rom[11823] = 8'hfa ;
            rom[11824] = 8'hd7 ;
            rom[11825] = 8'hc1 ;
            rom[11826] = 8'he0 ;
            rom[11827] = 8'h0c ;
            rom[11828] = 8'hf9 ;
            rom[11829] = 8'h0a ;
            rom[11830] = 8'h18 ;
            rom[11831] = 8'h01 ;
            rom[11832] = 8'heb ;
            rom[11833] = 8'he7 ;
            rom[11834] = 8'h27 ;
            rom[11835] = 8'hf0 ;
            rom[11836] = 8'h05 ;
            rom[11837] = 8'he8 ;
            rom[11838] = 8'h20 ;
            rom[11839] = 8'h16 ;
            rom[11840] = 8'hf1 ;
            rom[11841] = 8'h02 ;
            rom[11842] = 8'hda ;
            rom[11843] = 8'hf4 ;
            rom[11844] = 8'hee ;
            rom[11845] = 8'h0c ;
            rom[11846] = 8'he6 ;
            rom[11847] = 8'h1f ;
            rom[11848] = 8'hfe ;
            rom[11849] = 8'hed ;
            rom[11850] = 8'hfe ;
            rom[11851] = 8'h0a ;
            rom[11852] = 8'hbe ;
            rom[11853] = 8'h06 ;
            rom[11854] = 8'hf5 ;
            rom[11855] = 8'he9 ;
            rom[11856] = 8'h06 ;
            rom[11857] = 8'hf5 ;
            rom[11858] = 8'h41 ;
            rom[11859] = 8'hc0 ;
            rom[11860] = 8'h0a ;
            rom[11861] = 8'h07 ;
            rom[11862] = 8'h05 ;
            rom[11863] = 8'hfc ;
            rom[11864] = 8'hda ;
            rom[11865] = 8'hff ;
            rom[11866] = 8'hec ;
            rom[11867] = 8'h07 ;
            rom[11868] = 8'hce ;
            rom[11869] = 8'hd3 ;
            rom[11870] = 8'h1a ;
            rom[11871] = 8'h01 ;
            rom[11872] = 8'h11 ;
            rom[11873] = 8'h12 ;
            rom[11874] = 8'hd7 ;
            rom[11875] = 8'h26 ;
            rom[11876] = 8'hd1 ;
            rom[11877] = 8'he0 ;
            rom[11878] = 8'h05 ;
            rom[11879] = 8'he8 ;
            rom[11880] = 8'hfe ;
            rom[11881] = 8'h18 ;
            rom[11882] = 8'h01 ;
            rom[11883] = 8'hf7 ;
            rom[11884] = 8'hf8 ;
            rom[11885] = 8'heb ;
            rom[11886] = 8'h11 ;
            rom[11887] = 8'hdb ;
            rom[11888] = 8'hd1 ;
            rom[11889] = 8'h04 ;
            rom[11890] = 8'hff ;
            rom[11891] = 8'hf9 ;
            rom[11892] = 8'he5 ;
            rom[11893] = 8'h16 ;
            rom[11894] = 8'hed ;
            rom[11895] = 8'hfc ;
            rom[11896] = 8'h08 ;
            rom[11897] = 8'he8 ;
            rom[11898] = 8'h0c ;
            rom[11899] = 8'hf0 ;
            rom[11900] = 8'hf7 ;
            rom[11901] = 8'h0d ;
            rom[11902] = 8'hf4 ;
            rom[11903] = 8'hf5 ;
            rom[11904] = 8'h0d ;
            rom[11905] = 8'hf9 ;
            rom[11906] = 8'hdd ;
            rom[11907] = 8'h0a ;
            rom[11908] = 8'he8 ;
            rom[11909] = 8'he7 ;
            rom[11910] = 8'h08 ;
            rom[11911] = 8'heb ;
            rom[11912] = 8'h0d ;
            rom[11913] = 8'hfc ;
            rom[11914] = 8'he0 ;
            rom[11915] = 8'hf5 ;
            rom[11916] = 8'he0 ;
            rom[11917] = 8'hcc ;
            rom[11918] = 8'h0f ;
            rom[11919] = 8'h15 ;
            rom[11920] = 8'h0a ;
            rom[11921] = 8'hbb ;
            rom[11922] = 8'h0d ;
            rom[11923] = 8'hf2 ;
            rom[11924] = 8'hf1 ;
            rom[11925] = 8'h06 ;
            rom[11926] = 8'hfa ;
            rom[11927] = 8'hf8 ;
            rom[11928] = 8'hdd ;
            rom[11929] = 8'h19 ;
            rom[11930] = 8'h13 ;
            rom[11931] = 8'he5 ;
            rom[11932] = 8'h32 ;
            rom[11933] = 8'h00 ;
            rom[11934] = 8'h01 ;
            rom[11935] = 8'h0c ;
            rom[11936] = 8'h0f ;
            rom[11937] = 8'h12 ;
            rom[11938] = 8'hf3 ;
            rom[11939] = 8'hb8 ;
            rom[11940] = 8'hde ;
            rom[11941] = 8'hfc ;
            rom[11942] = 8'hf5 ;
            rom[11943] = 8'h11 ;
            rom[11944] = 8'hf0 ;
            rom[11945] = 8'hf0 ;
            rom[11946] = 8'hf8 ;
            rom[11947] = 8'h08 ;
            rom[11948] = 8'h18 ;
            rom[11949] = 8'h08 ;
            rom[11950] = 8'hf4 ;
            rom[11951] = 8'h24 ;
            rom[11952] = 8'hd9 ;
            rom[11953] = 8'hea ;
            rom[11954] = 8'he8 ;
            rom[11955] = 8'h0c ;
            rom[11956] = 8'hd8 ;
            rom[11957] = 8'hef ;
            rom[11958] = 8'hd6 ;
            rom[11959] = 8'hec ;
            rom[11960] = 8'h05 ;
            rom[11961] = 8'h09 ;
            rom[11962] = 8'hf4 ;
            rom[11963] = 8'hed ;
            rom[11964] = 8'he0 ;
            rom[11965] = 8'h17 ;
            rom[11966] = 8'hff ;
            rom[11967] = 8'hdf ;
            rom[11968] = 8'h0f ;
            rom[11969] = 8'hcf ;
            rom[11970] = 8'h17 ;
            rom[11971] = 8'he3 ;
            rom[11972] = 8'hed ;
            rom[11973] = 8'hef ;
            rom[11974] = 8'he0 ;
            rom[11975] = 8'he3 ;
            rom[11976] = 8'hfc ;
            rom[11977] = 8'hfb ;
            rom[11978] = 8'h0e ;
            rom[11979] = 8'heb ;
            rom[11980] = 8'h0e ;
            rom[11981] = 8'hfc ;
            rom[11982] = 8'hef ;
            rom[11983] = 8'h0e ;
            rom[11984] = 8'h1a ;
            rom[11985] = 8'h0c ;
            rom[11986] = 8'hf1 ;
            rom[11987] = 8'hf9 ;
            rom[11988] = 8'hf0 ;
            rom[11989] = 8'hfa ;
            rom[11990] = 8'hfb ;
            rom[11991] = 8'heb ;
            rom[11992] = 8'hfa ;
            rom[11993] = 8'h10 ;
            rom[11994] = 8'h0e ;
            rom[11995] = 8'h0a ;
            rom[11996] = 8'hdf ;
            rom[11997] = 8'hf4 ;
            rom[11998] = 8'hfe ;
            rom[11999] = 8'hfb ;
            rom[12000] = 8'h20 ;
            rom[12001] = 8'h01 ;
            rom[12002] = 8'hce ;
            rom[12003] = 8'he1 ;
            rom[12004] = 8'h02 ;
            rom[12005] = 8'hfd ;
            rom[12006] = 8'hf8 ;
            rom[12007] = 8'h03 ;
            rom[12008] = 8'h04 ;
            rom[12009] = 8'hf7 ;
            rom[12010] = 8'h0d ;
            rom[12011] = 8'hd1 ;
            rom[12012] = 8'h16 ;
            rom[12013] = 8'h15 ;
            rom[12014] = 8'h19 ;
            rom[12015] = 8'h13 ;
            rom[12016] = 8'h12 ;
            rom[12017] = 8'he8 ;
            rom[12018] = 8'h1d ;
            rom[12019] = 8'hef ;
            rom[12020] = 8'hf4 ;
            rom[12021] = 8'hed ;
            rom[12022] = 8'he9 ;
            rom[12023] = 8'hd9 ;
            rom[12024] = 8'he6 ;
            rom[12025] = 8'h1c ;
            rom[12026] = 8'h1b ;
            rom[12027] = 8'heb ;
            rom[12028] = 8'he3 ;
            rom[12029] = 8'he4 ;
            rom[12030] = 8'h06 ;
            rom[12031] = 8'hef ;
            rom[12032] = 8'hf1 ;
            rom[12033] = 8'hf3 ;
            rom[12034] = 8'hf7 ;
            rom[12035] = 8'h06 ;
            rom[12036] = 8'hf9 ;
            rom[12037] = 8'hff ;
            rom[12038] = 8'hf3 ;
            rom[12039] = 8'h02 ;
            rom[12040] = 8'h1d ;
            rom[12041] = 8'hfb ;
            rom[12042] = 8'hf4 ;
            rom[12043] = 8'hf9 ;
            rom[12044] = 8'hdd ;
            rom[12045] = 8'h01 ;
            rom[12046] = 8'heb ;
            rom[12047] = 8'hff ;
            rom[12048] = 8'he7 ;
            rom[12049] = 8'h03 ;
            rom[12050] = 8'h1c ;
            rom[12051] = 8'hea ;
            rom[12052] = 8'h2a ;
            rom[12053] = 8'h38 ;
            rom[12054] = 8'h10 ;
            rom[12055] = 8'hf2 ;
            rom[12056] = 8'h0c ;
            rom[12057] = 8'h1a ;
            rom[12058] = 8'hf9 ;
            rom[12059] = 8'hf9 ;
            rom[12060] = 8'hfc ;
            rom[12061] = 8'h15 ;
            rom[12062] = 8'heb ;
            rom[12063] = 8'h1f ;
            rom[12064] = 8'h1f ;
            rom[12065] = 8'h03 ;
            rom[12066] = 8'h15 ;
            rom[12067] = 8'hde ;
            rom[12068] = 8'h00 ;
            rom[12069] = 8'h03 ;
            rom[12070] = 8'h04 ;
            rom[12071] = 8'hfe ;
            rom[12072] = 8'h0b ;
            rom[12073] = 8'hd3 ;
            rom[12074] = 8'hf7 ;
            rom[12075] = 8'he3 ;
            rom[12076] = 8'h0d ;
            rom[12077] = 8'hda ;
            rom[12078] = 8'hfa ;
            rom[12079] = 8'hf9 ;
            rom[12080] = 8'hf2 ;
            rom[12081] = 8'h19 ;
            rom[12082] = 8'h04 ;
            rom[12083] = 8'hea ;
            rom[12084] = 8'hc9 ;
            rom[12085] = 8'hfb ;
            rom[12086] = 8'hff ;
            rom[12087] = 8'h0e ;
            rom[12088] = 8'h16 ;
            rom[12089] = 8'he9 ;
            rom[12090] = 8'h17 ;
            rom[12091] = 8'hec ;
            rom[12092] = 8'h14 ;
            rom[12093] = 8'h01 ;
            rom[12094] = 8'hd9 ;
            rom[12095] = 8'hed ;
            rom[12096] = 8'hf0 ;
            rom[12097] = 8'hdd ;
            rom[12098] = 8'h04 ;
            rom[12099] = 8'h04 ;
            rom[12100] = 8'h22 ;
            rom[12101] = 8'h2c ;
            rom[12102] = 8'h0e ;
            rom[12103] = 8'hf7 ;
            rom[12104] = 8'h22 ;
            rom[12105] = 8'hfc ;
            rom[12106] = 8'hec ;
            rom[12107] = 8'h29 ;
            rom[12108] = 8'h19 ;
            rom[12109] = 8'hdf ;
            rom[12110] = 8'hf1 ;
            rom[12111] = 8'he7 ;
            rom[12112] = 8'h13 ;
            rom[12113] = 8'hef ;
            rom[12114] = 8'hf7 ;
            rom[12115] = 8'hf4 ;
            rom[12116] = 8'hf9 ;
            rom[12117] = 8'hf4 ;
            rom[12118] = 8'hf5 ;
            rom[12119] = 8'he7 ;
            rom[12120] = 8'hff ;
            rom[12121] = 8'h0a ;
            rom[12122] = 8'h01 ;
            rom[12123] = 8'hd1 ;
            rom[12124] = 8'hef ;
            rom[12125] = 8'h03 ;
            rom[12126] = 8'hdb ;
            rom[12127] = 8'hc9 ;
            rom[12128] = 8'h07 ;
            rom[12129] = 8'h18 ;
            rom[12130] = 8'he7 ;
            rom[12131] = 8'hed ;
            rom[12132] = 8'hf5 ;
            rom[12133] = 8'h12 ;
            rom[12134] = 8'hfc ;
            rom[12135] = 8'he5 ;
            rom[12136] = 8'h12 ;
            rom[12137] = 8'h20 ;
            rom[12138] = 8'h09 ;
            rom[12139] = 8'h12 ;
            rom[12140] = 8'hfa ;
            rom[12141] = 8'h07 ;
            rom[12142] = 8'hf6 ;
            rom[12143] = 8'h0e ;
            rom[12144] = 8'hfa ;
            rom[12145] = 8'hff ;
            rom[12146] = 8'h21 ;
            rom[12147] = 8'h02 ;
            rom[12148] = 8'hf0 ;
            rom[12149] = 8'hfd ;
            rom[12150] = 8'he8 ;
            rom[12151] = 8'hea ;
            rom[12152] = 8'hc1 ;
            rom[12153] = 8'h15 ;
            rom[12154] = 8'hfb ;
            rom[12155] = 8'hef ;
            rom[12156] = 8'h1c ;
            rom[12157] = 8'h03 ;
            rom[12158] = 8'h30 ;
            rom[12159] = 8'h02 ;
            rom[12160] = 8'hf0 ;
            rom[12161] = 8'he8 ;
            rom[12162] = 8'h16 ;
            rom[12163] = 8'h0d ;
            rom[12164] = 8'hf0 ;
            rom[12165] = 8'hdf ;
            rom[12166] = 8'he9 ;
            rom[12167] = 8'h08 ;
            rom[12168] = 8'he7 ;
            rom[12169] = 8'hfa ;
            rom[12170] = 8'hf7 ;
            rom[12171] = 8'he8 ;
            rom[12172] = 8'hf3 ;
            rom[12173] = 8'hfd ;
            rom[12174] = 8'hf8 ;
            rom[12175] = 8'hc5 ;
            rom[12176] = 8'h0b ;
            rom[12177] = 8'hfa ;
            rom[12178] = 8'he4 ;
            rom[12179] = 8'h17 ;
            rom[12180] = 8'hd1 ;
            rom[12181] = 8'he1 ;
            rom[12182] = 8'h23 ;
            rom[12183] = 8'he7 ;
            rom[12184] = 8'hca ;
            rom[12185] = 8'heb ;
            rom[12186] = 8'h01 ;
            rom[12187] = 8'hd0 ;
            rom[12188] = 8'h15 ;
            rom[12189] = 8'hdf ;
            rom[12190] = 8'hd8 ;
            rom[12191] = 8'hfd ;
            rom[12192] = 8'hbd ;
            rom[12193] = 8'he2 ;
            rom[12194] = 8'he2 ;
            rom[12195] = 8'hf9 ;
            rom[12196] = 8'hf8 ;
            rom[12197] = 8'hee ;
            rom[12198] = 8'hfb ;
            rom[12199] = 8'hfb ;
            rom[12200] = 8'hf2 ;
            rom[12201] = 8'hea ;
            rom[12202] = 8'h02 ;
            rom[12203] = 8'hdf ;
            rom[12204] = 8'ha1 ;
            rom[12205] = 8'h0b ;
            rom[12206] = 8'hd1 ;
            rom[12207] = 8'he8 ;
            rom[12208] = 8'h12 ;
            rom[12209] = 8'hd2 ;
            rom[12210] = 8'h02 ;
            rom[12211] = 8'hf6 ;
            rom[12212] = 8'h04 ;
            rom[12213] = 8'h13 ;
            rom[12214] = 8'he7 ;
            rom[12215] = 8'hfd ;
            rom[12216] = 8'hd1 ;
            rom[12217] = 8'heb ;
            rom[12218] = 8'hca ;
            rom[12219] = 8'h32 ;
            rom[12220] = 8'hcf ;
            rom[12221] = 8'hfb ;
            rom[12222] = 8'hf0 ;
            rom[12223] = 8'hbf ;
            rom[12224] = 8'h00 ;
            rom[12225] = 8'hf3 ;
            rom[12226] = 8'hf4 ;
            rom[12227] = 8'hef ;
            rom[12228] = 8'h07 ;
            rom[12229] = 8'h05 ;
            rom[12230] = 8'hf8 ;
            rom[12231] = 8'h06 ;
            rom[12232] = 8'h12 ;
            rom[12233] = 8'he3 ;
            rom[12234] = 8'hfd ;
            rom[12235] = 8'h07 ;
            rom[12236] = 8'hed ;
            rom[12237] = 8'hf3 ;
            rom[12238] = 8'h14 ;
            rom[12239] = 8'h02 ;
            rom[12240] = 8'hec ;
            rom[12241] = 8'hf5 ;
            rom[12242] = 8'hf4 ;
            rom[12243] = 8'h16 ;
            rom[12244] = 8'h0f ;
            rom[12245] = 8'h0a ;
            rom[12246] = 8'hf0 ;
            rom[12247] = 8'h17 ;
            rom[12248] = 8'he9 ;
            rom[12249] = 8'he3 ;
            rom[12250] = 8'hee ;
            rom[12251] = 8'h15 ;
            rom[12252] = 8'hc7 ;
            rom[12253] = 8'hd8 ;
            rom[12254] = 8'hfd ;
            rom[12255] = 8'h05 ;
            rom[12256] = 8'hed ;
            rom[12257] = 8'hf2 ;
            rom[12258] = 8'hfd ;
            rom[12259] = 8'h00 ;
            rom[12260] = 8'hd8 ;
            rom[12261] = 8'hf8 ;
            rom[12262] = 8'he0 ;
            rom[12263] = 8'heb ;
            rom[12264] = 8'hdc ;
            rom[12265] = 8'hf8 ;
            rom[12266] = 8'he8 ;
            rom[12267] = 8'heb ;
            rom[12268] = 8'h1b ;
            rom[12269] = 8'h10 ;
            rom[12270] = 8'h20 ;
            rom[12271] = 8'h0e ;
            rom[12272] = 8'heb ;
            rom[12273] = 8'h1d ;
            rom[12274] = 8'hf3 ;
            rom[12275] = 8'hf6 ;
            rom[12276] = 8'h9d ;
            rom[12277] = 8'h1a ;
            rom[12278] = 8'hed ;
            rom[12279] = 8'h0c ;
            rom[12280] = 8'hf5 ;
            rom[12281] = 8'h03 ;
            rom[12282] = 8'he2 ;
            rom[12283] = 8'hfc ;
            rom[12284] = 8'heb ;
            rom[12285] = 8'he3 ;
            rom[12286] = 8'he6 ;
            rom[12287] = 8'hd8 ;
            rom[12288] = 8'he7 ;
            rom[12289] = 8'h0a ;
            rom[12290] = 8'he6 ;
            rom[12291] = 8'h13 ;
            rom[12292] = 8'h08 ;
            rom[12293] = 8'h1c ;
            rom[12294] = 8'he2 ;
            rom[12295] = 8'hef ;
            rom[12296] = 8'h14 ;
            rom[12297] = 8'hea ;
            rom[12298] = 8'h06 ;
            rom[12299] = 8'hfb ;
            rom[12300] = 8'hda ;
            rom[12301] = 8'h1d ;
            rom[12302] = 8'h0c ;
            rom[12303] = 8'h01 ;
            rom[12304] = 8'hea ;
            rom[12305] = 8'hf2 ;
            rom[12306] = 8'hfb ;
            rom[12307] = 8'h01 ;
            rom[12308] = 8'h02 ;
            rom[12309] = 8'hf6 ;
            rom[12310] = 8'h1c ;
            rom[12311] = 8'he2 ;
            rom[12312] = 8'h16 ;
            rom[12313] = 8'h32 ;
            rom[12314] = 8'h02 ;
            rom[12315] = 8'hee ;
            rom[12316] = 8'h0f ;
            rom[12317] = 8'h0a ;
            rom[12318] = 8'h04 ;
            rom[12319] = 8'hf3 ;
            rom[12320] = 8'h1b ;
            rom[12321] = 8'h17 ;
            rom[12322] = 8'he4 ;
            rom[12323] = 8'hc9 ;
            rom[12324] = 8'hd8 ;
            rom[12325] = 8'hca ;
            rom[12326] = 8'hfd ;
            rom[12327] = 8'h08 ;
            rom[12328] = 8'h0a ;
            rom[12329] = 8'hcb ;
            rom[12330] = 8'hf4 ;
            rom[12331] = 8'heb ;
            rom[12332] = 8'h14 ;
            rom[12333] = 8'h00 ;
            rom[12334] = 8'he1 ;
            rom[12335] = 8'hec ;
            rom[12336] = 8'he7 ;
            rom[12337] = 8'h11 ;
            rom[12338] = 8'hd7 ;
            rom[12339] = 8'hd6 ;
            rom[12340] = 8'hca ;
            rom[12341] = 8'hce ;
            rom[12342] = 8'h15 ;
            rom[12343] = 8'h0e ;
            rom[12344] = 8'hff ;
            rom[12345] = 8'hfc ;
            rom[12346] = 8'h00 ;
            rom[12347] = 8'he5 ;
            rom[12348] = 8'h13 ;
            rom[12349] = 8'h0f ;
            rom[12350] = 8'hf1 ;
            rom[12351] = 8'h06 ;
            rom[12352] = 8'h12 ;
            rom[12353] = 8'heb ;
            rom[12354] = 8'h32 ;
            rom[12355] = 8'hee ;
            rom[12356] = 8'h08 ;
            rom[12357] = 8'h26 ;
            rom[12358] = 8'he1 ;
            rom[12359] = 8'hcb ;
            rom[12360] = 8'h03 ;
            rom[12361] = 8'h0a ;
            rom[12362] = 8'hde ;
            rom[12363] = 8'he1 ;
            rom[12364] = 8'h05 ;
            rom[12365] = 8'he2 ;
            rom[12366] = 8'he8 ;
            rom[12367] = 8'h16 ;
            rom[12368] = 8'h1a ;
            rom[12369] = 8'hdb ;
            rom[12370] = 8'h26 ;
            rom[12371] = 8'hf0 ;
            rom[12372] = 8'hf1 ;
            rom[12373] = 8'h1d ;
            rom[12374] = 8'he1 ;
            rom[12375] = 8'hf4 ;
            rom[12376] = 8'he7 ;
            rom[12377] = 8'he1 ;
            rom[12378] = 8'hec ;
            rom[12379] = 8'hed ;
            rom[12380] = 8'h01 ;
            rom[12381] = 8'h0f ;
            rom[12382] = 8'hf6 ;
            rom[12383] = 8'hd1 ;
            rom[12384] = 8'h0c ;
            rom[12385] = 8'h0e ;
            rom[12386] = 8'h02 ;
            rom[12387] = 8'h0d ;
            rom[12388] = 8'h1c ;
            rom[12389] = 8'hfa ;
            rom[12390] = 8'h07 ;
            rom[12391] = 8'hf5 ;
            rom[12392] = 8'hde ;
            rom[12393] = 8'hf0 ;
            rom[12394] = 8'h21 ;
            rom[12395] = 8'hf7 ;
            rom[12396] = 8'h22 ;
            rom[12397] = 8'h1d ;
            rom[12398] = 8'h02 ;
            rom[12399] = 8'he1 ;
            rom[12400] = 8'h0e ;
            rom[12401] = 8'h07 ;
            rom[12402] = 8'h2e ;
            rom[12403] = 8'hfb ;
            rom[12404] = 8'h09 ;
            rom[12405] = 8'hc7 ;
            rom[12406] = 8'heb ;
            rom[12407] = 8'hcc ;
            rom[12408] = 8'he0 ;
            rom[12409] = 8'h14 ;
            rom[12410] = 8'he7 ;
            rom[12411] = 8'h0d ;
            rom[12412] = 8'hcc ;
            rom[12413] = 8'h14 ;
            rom[12414] = 8'h09 ;
            rom[12415] = 8'h0d ;
            rom[12416] = 8'h1b ;
            rom[12417] = 8'hd2 ;
            rom[12418] = 8'h10 ;
            rom[12419] = 8'h1c ;
            rom[12420] = 8'h00 ;
            rom[12421] = 8'hf5 ;
            rom[12422] = 8'hd6 ;
            rom[12423] = 8'hd9 ;
            rom[12424] = 8'hf4 ;
            rom[12425] = 8'h1a ;
            rom[12426] = 8'h01 ;
            rom[12427] = 8'hf3 ;
            rom[12428] = 8'he7 ;
            rom[12429] = 8'he9 ;
            rom[12430] = 8'h08 ;
            rom[12431] = 8'hf8 ;
            rom[12432] = 8'hdc ;
            rom[12433] = 8'h06 ;
            rom[12434] = 8'h06 ;
            rom[12435] = 8'hdb ;
            rom[12436] = 8'hef ;
            rom[12437] = 8'hdc ;
            rom[12438] = 8'h09 ;
            rom[12439] = 8'hfa ;
            rom[12440] = 8'h01 ;
            rom[12441] = 8'he0 ;
            rom[12442] = 8'h13 ;
            rom[12443] = 8'hd8 ;
            rom[12444] = 8'hd5 ;
            rom[12445] = 8'h25 ;
            rom[12446] = 8'he1 ;
            rom[12447] = 8'h1a ;
            rom[12448] = 8'he5 ;
            rom[12449] = 8'h09 ;
            rom[12450] = 8'hc8 ;
            rom[12451] = 8'hec ;
            rom[12452] = 8'hfd ;
            rom[12453] = 8'hd8 ;
            rom[12454] = 8'hd4 ;
            rom[12455] = 8'h00 ;
            rom[12456] = 8'hf4 ;
            rom[12457] = 8'hdb ;
            rom[12458] = 8'h01 ;
            rom[12459] = 8'hf0 ;
            rom[12460] = 8'h14 ;
            rom[12461] = 8'h2c ;
            rom[12462] = 8'h03 ;
            rom[12463] = 8'hd8 ;
            rom[12464] = 8'hc8 ;
            rom[12465] = 8'he6 ;
            rom[12466] = 8'hfb ;
            rom[12467] = 8'hef ;
            rom[12468] = 8'h1b ;
            rom[12469] = 8'h09 ;
            rom[12470] = 8'h0d ;
            rom[12471] = 8'hd6 ;
            rom[12472] = 8'h12 ;
            rom[12473] = 8'h17 ;
            rom[12474] = 8'h1f ;
            rom[12475] = 8'he3 ;
            rom[12476] = 8'hfc ;
            rom[12477] = 8'hd1 ;
            rom[12478] = 8'h06 ;
            rom[12479] = 8'hec ;
            rom[12480] = 8'hd3 ;
            rom[12481] = 8'h11 ;
            rom[12482] = 8'h19 ;
            rom[12483] = 8'h1d ;
            rom[12484] = 8'hf9 ;
            rom[12485] = 8'hf9 ;
            rom[12486] = 8'hd6 ;
            rom[12487] = 8'h0e ;
            rom[12488] = 8'h0c ;
            rom[12489] = 8'he6 ;
            rom[12490] = 8'h12 ;
            rom[12491] = 8'hed ;
            rom[12492] = 8'hf8 ;
            rom[12493] = 8'h11 ;
            rom[12494] = 8'h07 ;
            rom[12495] = 8'h02 ;
            rom[12496] = 8'hfe ;
            rom[12497] = 8'h02 ;
            rom[12498] = 8'hf1 ;
            rom[12499] = 8'hdb ;
            rom[12500] = 8'hf6 ;
            rom[12501] = 8'hda ;
            rom[12502] = 8'he6 ;
            rom[12503] = 8'hf7 ;
            rom[12504] = 8'h14 ;
            rom[12505] = 8'hec ;
            rom[12506] = 8'hff ;
            rom[12507] = 8'h05 ;
            rom[12508] = 8'h08 ;
            rom[12509] = 8'hf0 ;
            rom[12510] = 8'h1d ;
            rom[12511] = 8'hf6 ;
            rom[12512] = 8'h02 ;
            rom[12513] = 8'hf4 ;
            rom[12514] = 8'hf6 ;
            rom[12515] = 8'heb ;
            rom[12516] = 8'he9 ;
            rom[12517] = 8'he7 ;
            rom[12518] = 8'h0b ;
            rom[12519] = 8'hfb ;
            rom[12520] = 8'hee ;
            rom[12521] = 8'h0e ;
            rom[12522] = 8'he8 ;
            rom[12523] = 8'h04 ;
            rom[12524] = 8'hf0 ;
            rom[12525] = 8'h0d ;
            rom[12526] = 8'h0e ;
            rom[12527] = 8'hf9 ;
            rom[12528] = 8'hec ;
            rom[12529] = 8'hf6 ;
            rom[12530] = 8'h03 ;
            rom[12531] = 8'h01 ;
            rom[12532] = 8'hfc ;
            rom[12533] = 8'hf8 ;
            rom[12534] = 8'h0d ;
            rom[12535] = 8'hf8 ;
            rom[12536] = 8'h15 ;
            rom[12537] = 8'h0b ;
            rom[12538] = 8'h10 ;
            rom[12539] = 8'hda ;
            rom[12540] = 8'hf2 ;
            rom[12541] = 8'he8 ;
            rom[12542] = 8'haf ;
            rom[12543] = 8'hf9 ;
            rom[12544] = 8'h19 ;
            rom[12545] = 8'he8 ;
            rom[12546] = 8'hfb ;
            rom[12547] = 8'h03 ;
            rom[12548] = 8'h01 ;
            rom[12549] = 8'h03 ;
            rom[12550] = 8'hcb ;
            rom[12551] = 8'hde ;
            rom[12552] = 8'h01 ;
            rom[12553] = 8'h05 ;
            rom[12554] = 8'hfc ;
            rom[12555] = 8'hea ;
            rom[12556] = 8'hde ;
            rom[12557] = 8'hef ;
            rom[12558] = 8'h0a ;
            rom[12559] = 8'he2 ;
            rom[12560] = 8'h0f ;
            rom[12561] = 8'h08 ;
            rom[12562] = 8'h0d ;
            rom[12563] = 8'h01 ;
            rom[12564] = 8'hfd ;
            rom[12565] = 8'hd9 ;
            rom[12566] = 8'hf4 ;
            rom[12567] = 8'hf3 ;
            rom[12568] = 8'h21 ;
            rom[12569] = 8'he9 ;
            rom[12570] = 8'hf5 ;
            rom[12571] = 8'he5 ;
            rom[12572] = 8'hff ;
            rom[12573] = 8'h13 ;
            rom[12574] = 8'h08 ;
            rom[12575] = 8'h02 ;
            rom[12576] = 8'h0d ;
            rom[12577] = 8'h03 ;
            rom[12578] = 8'h07 ;
            rom[12579] = 8'hdd ;
            rom[12580] = 8'h06 ;
            rom[12581] = 8'hf8 ;
            rom[12582] = 8'he7 ;
            rom[12583] = 8'he9 ;
            rom[12584] = 8'hf9 ;
            rom[12585] = 8'h1f ;
            rom[12586] = 8'hf3 ;
            rom[12587] = 8'hf2 ;
            rom[12588] = 8'h0c ;
            rom[12589] = 8'h00 ;
            rom[12590] = 8'h19 ;
            rom[12591] = 8'hcf ;
            rom[12592] = 8'hf8 ;
            rom[12593] = 8'hff ;
            rom[12594] = 8'hf4 ;
            rom[12595] = 8'h03 ;
            rom[12596] = 8'h09 ;
            rom[12597] = 8'hf7 ;
            rom[12598] = 8'hec ;
            rom[12599] = 8'h07 ;
            rom[12600] = 8'h10 ;
            rom[12601] = 8'h03 ;
            rom[12602] = 8'hff ;
            rom[12603] = 8'h12 ;
            rom[12604] = 8'h19 ;
            rom[12605] = 8'hc6 ;
            rom[12606] = 8'hf3 ;
            rom[12607] = 8'hfb ;
            rom[12608] = 8'hf3 ;
            rom[12609] = 8'h05 ;
            rom[12610] = 8'h19 ;
            rom[12611] = 8'hee ;
            rom[12612] = 8'hec ;
            rom[12613] = 8'hff ;
            rom[12614] = 8'hfe ;
            rom[12615] = 8'he0 ;
            rom[12616] = 8'h0e ;
            rom[12617] = 8'h03 ;
            rom[12618] = 8'hf3 ;
            rom[12619] = 8'h0a ;
            rom[12620] = 8'hfe ;
            rom[12621] = 8'h19 ;
            rom[12622] = 8'hfa ;
            rom[12623] = 8'hd7 ;
            rom[12624] = 8'hd5 ;
            rom[12625] = 8'h14 ;
            rom[12626] = 8'h00 ;
            rom[12627] = 8'he6 ;
            rom[12628] = 8'h03 ;
            rom[12629] = 8'h23 ;
            rom[12630] = 8'hc5 ;
            rom[12631] = 8'hfa ;
            rom[12632] = 8'he0 ;
            rom[12633] = 8'hea ;
            rom[12634] = 8'hd0 ;
            rom[12635] = 8'h03 ;
            rom[12636] = 8'hd3 ;
            rom[12637] = 8'h05 ;
            rom[12638] = 8'hd9 ;
            rom[12639] = 8'h02 ;
            rom[12640] = 8'he9 ;
            rom[12641] = 8'hd7 ;
            rom[12642] = 8'h1b ;
            rom[12643] = 8'h1f ;
            rom[12644] = 8'h07 ;
            rom[12645] = 8'h0f ;
            rom[12646] = 8'h00 ;
            rom[12647] = 8'hf5 ;
            rom[12648] = 8'hf1 ;
            rom[12649] = 8'hf8 ;
            rom[12650] = 8'h33 ;
            rom[12651] = 8'hff ;
            rom[12652] = 8'h1f ;
            rom[12653] = 8'hf7 ;
            rom[12654] = 8'h13 ;
            rom[12655] = 8'hed ;
            rom[12656] = 8'hd8 ;
            rom[12657] = 8'he4 ;
            rom[12658] = 8'h30 ;
            rom[12659] = 8'he6 ;
            rom[12660] = 8'h28 ;
            rom[12661] = 8'h08 ;
            rom[12662] = 8'hdc ;
            rom[12663] = 8'hfa ;
            rom[12664] = 8'hea ;
            rom[12665] = 8'hd1 ;
            rom[12666] = 8'he9 ;
            rom[12667] = 8'h15 ;
            rom[12668] = 8'h0b ;
            rom[12669] = 8'hfb ;
            rom[12670] = 8'hfd ;
            rom[12671] = 8'hcb ;
            rom[12672] = 8'h28 ;
            rom[12673] = 8'hc0 ;
            rom[12674] = 8'h29 ;
            rom[12675] = 8'h2d ;
            rom[12676] = 8'he4 ;
            rom[12677] = 8'hf7 ;
            rom[12678] = 8'h06 ;
            rom[12679] = 8'hf7 ;
            rom[12680] = 8'hef ;
            rom[12681] = 8'he6 ;
            rom[12682] = 8'h07 ;
            rom[12683] = 8'h04 ;
            rom[12684] = 8'h13 ;
            rom[12685] = 8'h12 ;
            rom[12686] = 8'hfa ;
            rom[12687] = 8'h07 ;
            rom[12688] = 8'hd9 ;
            rom[12689] = 8'hf3 ;
            rom[12690] = 8'h04 ;
            rom[12691] = 8'h1b ;
            rom[12692] = 8'h0e ;
            rom[12693] = 8'hc8 ;
            rom[12694] = 8'hf3 ;
            rom[12695] = 8'hd9 ;
            rom[12696] = 8'h17 ;
            rom[12697] = 8'hce ;
            rom[12698] = 8'h2c ;
            rom[12699] = 8'hd0 ;
            rom[12700] = 8'hf9 ;
            rom[12701] = 8'hf4 ;
            rom[12702] = 8'hee ;
            rom[12703] = 8'h0c ;
            rom[12704] = 8'heb ;
            rom[12705] = 8'hfe ;
            rom[12706] = 8'hec ;
            rom[12707] = 8'h03 ;
            rom[12708] = 8'h1c ;
            rom[12709] = 8'hed ;
            rom[12710] = 8'h07 ;
            rom[12711] = 8'he8 ;
            rom[12712] = 8'h16 ;
            rom[12713] = 8'he3 ;
            rom[12714] = 8'hfa ;
            rom[12715] = 8'hfd ;
            rom[12716] = 8'hf1 ;
            rom[12717] = 8'h0c ;
            rom[12718] = 8'hf7 ;
            rom[12719] = 8'hdc ;
            rom[12720] = 8'hd8 ;
            rom[12721] = 8'hf7 ;
            rom[12722] = 8'hf7 ;
            rom[12723] = 8'h00 ;
            rom[12724] = 8'h15 ;
            rom[12725] = 8'hf0 ;
            rom[12726] = 8'hc2 ;
            rom[12727] = 8'h01 ;
            rom[12728] = 8'h11 ;
            rom[12729] = 8'h26 ;
            rom[12730] = 8'h03 ;
            rom[12731] = 8'hf0 ;
            rom[12732] = 8'h04 ;
            rom[12733] = 8'h12 ;
            rom[12734] = 8'he8 ;
            rom[12735] = 8'hd5 ;
            rom[12736] = 8'hd4 ;
            rom[12737] = 8'h19 ;
            rom[12738] = 8'hfb ;
            rom[12739] = 8'hee ;
            rom[12740] = 8'h07 ;
            rom[12741] = 8'h19 ;
            rom[12742] = 8'hdb ;
            rom[12743] = 8'h01 ;
            rom[12744] = 8'h0b ;
            rom[12745] = 8'h0d ;
            rom[12746] = 8'hcf ;
            rom[12747] = 8'hfd ;
            rom[12748] = 8'he5 ;
            rom[12749] = 8'h34 ;
            rom[12750] = 8'h1a ;
            rom[12751] = 8'h0a ;
            rom[12752] = 8'h00 ;
            rom[12753] = 8'h1c ;
            rom[12754] = 8'heb ;
            rom[12755] = 8'he4 ;
            rom[12756] = 8'hf1 ;
            rom[12757] = 8'hdf ;
            rom[12758] = 8'hfd ;
            rom[12759] = 8'he8 ;
            rom[12760] = 8'hfa ;
            rom[12761] = 8'hed ;
            rom[12762] = 8'h1b ;
            rom[12763] = 8'h11 ;
            rom[12764] = 8'h22 ;
            rom[12765] = 8'hfd ;
            rom[12766] = 8'h13 ;
            rom[12767] = 8'hf6 ;
            rom[12768] = 8'heb ;
            rom[12769] = 8'h08 ;
            rom[12770] = 8'h01 ;
            rom[12771] = 8'h0f ;
            rom[12772] = 8'he7 ;
            rom[12773] = 8'h07 ;
            rom[12774] = 8'hf7 ;
            rom[12775] = 8'hdf ;
            rom[12776] = 8'hed ;
            rom[12777] = 8'hfa ;
            rom[12778] = 8'h04 ;
            rom[12779] = 8'hfd ;
            rom[12780] = 8'hfe ;
            rom[12781] = 8'h0c ;
            rom[12782] = 8'h0a ;
            rom[12783] = 8'he5 ;
            rom[12784] = 8'hf1 ;
            rom[12785] = 8'he0 ;
            rom[12786] = 8'h1f ;
            rom[12787] = 8'h0e ;
            rom[12788] = 8'hfa ;
            rom[12789] = 8'hfd ;
            rom[12790] = 8'he5 ;
            rom[12791] = 8'he6 ;
            rom[12792] = 8'hfa ;
            rom[12793] = 8'he2 ;
            rom[12794] = 8'hf1 ;
            rom[12795] = 8'hf7 ;
            rom[12796] = 8'hdc ;
            rom[12797] = 8'hed ;
            rom[12798] = 8'he6 ;
            rom[12799] = 8'h10 ;
            rom[12800] = 8'hea ;
            rom[12801] = 8'hfe ;
            rom[12802] = 8'h0f ;
            rom[12803] = 8'hf5 ;
            rom[12804] = 8'hf5 ;
            rom[12805] = 8'heb ;
            rom[12806] = 8'h11 ;
            rom[12807] = 8'h14 ;
            rom[12808] = 8'hda ;
            rom[12809] = 8'hf5 ;
            rom[12810] = 8'hf1 ;
            rom[12811] = 8'hfd ;
            rom[12812] = 8'h25 ;
            rom[12813] = 8'h03 ;
            rom[12814] = 8'hd8 ;
            rom[12815] = 8'hf1 ;
            rom[12816] = 8'he4 ;
            rom[12817] = 8'hff ;
            rom[12818] = 8'hf3 ;
            rom[12819] = 8'hc9 ;
            rom[12820] = 8'h0a ;
            rom[12821] = 8'h07 ;
            rom[12822] = 8'h06 ;
            rom[12823] = 8'hfe ;
            rom[12824] = 8'h12 ;
            rom[12825] = 8'hf7 ;
            rom[12826] = 8'hdb ;
            rom[12827] = 8'h10 ;
            rom[12828] = 8'hfd ;
            rom[12829] = 8'h20 ;
            rom[12830] = 8'h04 ;
            rom[12831] = 8'h1b ;
            rom[12832] = 8'h22 ;
            rom[12833] = 8'hda ;
            rom[12834] = 8'hf9 ;
            rom[12835] = 8'hfd ;
            rom[12836] = 8'hef ;
            rom[12837] = 8'hda ;
            rom[12838] = 8'h10 ;
            rom[12839] = 8'he0 ;
            rom[12840] = 8'h1c ;
            rom[12841] = 8'hd8 ;
            rom[12842] = 8'hf1 ;
            rom[12843] = 8'he9 ;
            rom[12844] = 8'h09 ;
            rom[12845] = 8'hff ;
            rom[12846] = 8'hc3 ;
            rom[12847] = 8'h0d ;
            rom[12848] = 8'h23 ;
            rom[12849] = 8'h02 ;
            rom[12850] = 8'h03 ;
            rom[12851] = 8'h09 ;
            rom[12852] = 8'h12 ;
            rom[12853] = 8'h0d ;
            rom[12854] = 8'he2 ;
            rom[12855] = 8'hda ;
            rom[12856] = 8'hf6 ;
            rom[12857] = 8'hf8 ;
            rom[12858] = 8'hdf ;
            rom[12859] = 8'h1a ;
            rom[12860] = 8'hf7 ;
            rom[12861] = 8'h05 ;
            rom[12862] = 8'hdd ;
            rom[12863] = 8'h07 ;
            rom[12864] = 8'h03 ;
            rom[12865] = 8'hfc ;
            rom[12866] = 8'hf2 ;
            rom[12867] = 8'he5 ;
            rom[12868] = 8'h04 ;
            rom[12869] = 8'he2 ;
            rom[12870] = 8'h0c ;
            rom[12871] = 8'h12 ;
            rom[12872] = 8'hea ;
            rom[12873] = 8'hf9 ;
            rom[12874] = 8'hf0 ;
            rom[12875] = 8'he9 ;
            rom[12876] = 8'hdc ;
            rom[12877] = 8'had ;
            rom[12878] = 8'hec ;
            rom[12879] = 8'h04 ;
            rom[12880] = 8'he8 ;
            rom[12881] = 8'hfe ;
            rom[12882] = 8'hee ;
            rom[12883] = 8'hfb ;
            rom[12884] = 8'hd4 ;
            rom[12885] = 8'hf5 ;
            rom[12886] = 8'hf9 ;
            rom[12887] = 8'hef ;
            rom[12888] = 8'he5 ;
            rom[12889] = 8'h06 ;
            rom[12890] = 8'hfa ;
            rom[12891] = 8'hef ;
            rom[12892] = 8'hf1 ;
            rom[12893] = 8'h00 ;
            rom[12894] = 8'he3 ;
            rom[12895] = 8'hfd ;
            rom[12896] = 8'he6 ;
            rom[12897] = 8'h01 ;
            rom[12898] = 8'he0 ;
            rom[12899] = 8'h02 ;
            rom[12900] = 8'h01 ;
            rom[12901] = 8'h10 ;
            rom[12902] = 8'h0f ;
            rom[12903] = 8'he6 ;
            rom[12904] = 8'he9 ;
            rom[12905] = 8'h09 ;
            rom[12906] = 8'hfc ;
            rom[12907] = 8'h05 ;
            rom[12908] = 8'he0 ;
            rom[12909] = 8'hf1 ;
            rom[12910] = 8'hf5 ;
            rom[12911] = 8'h1d ;
            rom[12912] = 8'h07 ;
            rom[12913] = 8'hf3 ;
            rom[12914] = 8'hf1 ;
            rom[12915] = 8'hfd ;
            rom[12916] = 8'hec ;
            rom[12917] = 8'h1e ;
            rom[12918] = 8'h02 ;
            rom[12919] = 8'hf2 ;
            rom[12920] = 8'hd6 ;
            rom[12921] = 8'h0a ;
            rom[12922] = 8'h03 ;
            rom[12923] = 8'hf6 ;
            rom[12924] = 8'hfb ;
            rom[12925] = 8'he7 ;
            rom[12926] = 8'hc6 ;
            rom[12927] = 8'h11 ;
            rom[12928] = 8'hd1 ;
            rom[12929] = 8'h0f ;
            rom[12930] = 8'h0b ;
            rom[12931] = 8'hf7 ;
            rom[12932] = 8'h18 ;
            rom[12933] = 8'h15 ;
            rom[12934] = 8'hfa ;
            rom[12935] = 8'hf4 ;
            rom[12936] = 8'hf8 ;
            rom[12937] = 8'he7 ;
            rom[12938] = 8'hf0 ;
            rom[12939] = 8'hfe ;
            rom[12940] = 8'h0c ;
            rom[12941] = 8'h17 ;
            rom[12942] = 8'hf5 ;
            rom[12943] = 8'h0c ;
            rom[12944] = 8'hfe ;
            rom[12945] = 8'hf7 ;
            rom[12946] = 8'hc2 ;
            rom[12947] = 8'hbc ;
            rom[12948] = 8'hfc ;
            rom[12949] = 8'hf7 ;
            rom[12950] = 8'h10 ;
            rom[12951] = 8'h14 ;
            rom[12952] = 8'h24 ;
            rom[12953] = 8'hf6 ;
            rom[12954] = 8'h12 ;
            rom[12955] = 8'h1f ;
            rom[12956] = 8'hff ;
            rom[12957] = 8'hf3 ;
            rom[12958] = 8'hed ;
            rom[12959] = 8'ha9 ;
            rom[12960] = 8'h13 ;
            rom[12961] = 8'he5 ;
            rom[12962] = 8'h22 ;
            rom[12963] = 8'hf5 ;
            rom[12964] = 8'hf6 ;
            rom[12965] = 8'h16 ;
            rom[12966] = 8'h0c ;
            rom[12967] = 8'hfe ;
            rom[12968] = 8'hf8 ;
            rom[12969] = 8'hed ;
            rom[12970] = 8'hd7 ;
            rom[12971] = 8'hf5 ;
            rom[12972] = 8'h0a ;
            rom[12973] = 8'h0e ;
            rom[12974] = 8'h36 ;
            rom[12975] = 8'h0b ;
            rom[12976] = 8'he5 ;
            rom[12977] = 8'h23 ;
            rom[12978] = 8'h01 ;
            rom[12979] = 8'he6 ;
            rom[12980] = 8'hee ;
            rom[12981] = 8'hf4 ;
            rom[12982] = 8'h06 ;
            rom[12983] = 8'hee ;
            rom[12984] = 8'h35 ;
            rom[12985] = 8'hf7 ;
            rom[12986] = 8'hf0 ;
            rom[12987] = 8'he0 ;
            rom[12988] = 8'hf0 ;
            rom[12989] = 8'he1 ;
            rom[12990] = 8'he1 ;
            rom[12991] = 8'hfc ;
            rom[12992] = 8'h02 ;
            rom[12993] = 8'hfa ;
            rom[12994] = 8'he3 ;
            rom[12995] = 8'h04 ;
            rom[12996] = 8'hed ;
            rom[12997] = 8'hee ;
            rom[12998] = 8'h11 ;
            rom[12999] = 8'h12 ;
            rom[13000] = 8'hc6 ;
            rom[13001] = 8'hdd ;
            rom[13002] = 8'h09 ;
            rom[13003] = 8'h1d ;
            rom[13004] = 8'hda ;
            rom[13005] = 8'he9 ;
            rom[13006] = 8'hc6 ;
            rom[13007] = 8'h04 ;
            rom[13008] = 8'h03 ;
            rom[13009] = 8'h07 ;
            rom[13010] = 8'h15 ;
            rom[13011] = 8'h0e ;
            rom[13012] = 8'h0d ;
            rom[13013] = 8'h09 ;
            rom[13014] = 8'hf4 ;
            rom[13015] = 8'hcb ;
            rom[13016] = 8'h23 ;
            rom[13017] = 8'h05 ;
            rom[13018] = 8'h01 ;
            rom[13019] = 8'h01 ;
            rom[13020] = 8'h16 ;
            rom[13021] = 8'h37 ;
            rom[13022] = 8'hf1 ;
            rom[13023] = 8'hf6 ;
            rom[13024] = 8'hd5 ;
            rom[13025] = 8'hed ;
            rom[13026] = 8'h07 ;
            rom[13027] = 8'hd6 ;
            rom[13028] = 8'h09 ;
            rom[13029] = 8'hf2 ;
            rom[13030] = 8'h0d ;
            rom[13031] = 8'h10 ;
            rom[13032] = 8'h17 ;
            rom[13033] = 8'hed ;
            rom[13034] = 8'hff ;
            rom[13035] = 8'h07 ;
            rom[13036] = 8'h06 ;
            rom[13037] = 8'hf5 ;
            rom[13038] = 8'hdc ;
            rom[13039] = 8'h18 ;
            rom[13040] = 8'hff ;
            rom[13041] = 8'h04 ;
            rom[13042] = 8'h29 ;
            rom[13043] = 8'h16 ;
            rom[13044] = 8'hfe ;
            rom[13045] = 8'h0f ;
            rom[13046] = 8'hf5 ;
            rom[13047] = 8'h0c ;
            rom[13048] = 8'hd1 ;
            rom[13049] = 8'he9 ;
            rom[13050] = 8'hfc ;
            rom[13051] = 8'he0 ;
            rom[13052] = 8'h0e ;
            rom[13053] = 8'h0f ;
            rom[13054] = 8'h11 ;
            rom[13055] = 8'hfb ;
            rom[13056] = 8'hf9 ;
            rom[13057] = 8'hf8 ;
            rom[13058] = 8'he5 ;
            rom[13059] = 8'h05 ;
            rom[13060] = 8'h10 ;
            rom[13061] = 8'h02 ;
            rom[13062] = 8'hf3 ;
            rom[13063] = 8'h0e ;
            rom[13064] = 8'h1e ;
            rom[13065] = 8'hf2 ;
            rom[13066] = 8'h02 ;
            rom[13067] = 8'h06 ;
            rom[13068] = 8'h09 ;
            rom[13069] = 8'hc9 ;
            rom[13070] = 8'h09 ;
            rom[13071] = 8'h0b ;
            rom[13072] = 8'heb ;
            rom[13073] = 8'hf0 ;
            rom[13074] = 8'h19 ;
            rom[13075] = 8'h1c ;
            rom[13076] = 8'hed ;
            rom[13077] = 8'hd5 ;
            rom[13078] = 8'hf9 ;
            rom[13079] = 8'h10 ;
            rom[13080] = 8'h21 ;
            rom[13081] = 8'h12 ;
            rom[13082] = 8'h1a ;
            rom[13083] = 8'hfe ;
            rom[13084] = 8'hf7 ;
            rom[13085] = 8'h0f ;
            rom[13086] = 8'hed ;
            rom[13087] = 8'hed ;
            rom[13088] = 8'h00 ;
            rom[13089] = 8'hb6 ;
            rom[13090] = 8'he1 ;
            rom[13091] = 8'hfa ;
            rom[13092] = 8'h0a ;
            rom[13093] = 8'hf3 ;
            rom[13094] = 8'hf1 ;
            rom[13095] = 8'h04 ;
            rom[13096] = 8'h2a ;
            rom[13097] = 8'he1 ;
            rom[13098] = 8'he6 ;
            rom[13099] = 8'hdd ;
            rom[13100] = 8'h08 ;
            rom[13101] = 8'h01 ;
            rom[13102] = 8'he7 ;
            rom[13103] = 8'hde ;
            rom[13104] = 8'hc9 ;
            rom[13105] = 8'h03 ;
            rom[13106] = 8'hf1 ;
            rom[13107] = 8'hea ;
            rom[13108] = 8'h01 ;
            rom[13109] = 8'hf4 ;
            rom[13110] = 8'h06 ;
            rom[13111] = 8'hf5 ;
            rom[13112] = 8'he0 ;
            rom[13113] = 8'h1a ;
            rom[13114] = 8'h14 ;
            rom[13115] = 8'h10 ;
            rom[13116] = 8'h12 ;
            rom[13117] = 8'hf9 ;
            rom[13118] = 8'h18 ;
            rom[13119] = 8'hf6 ;
            rom[13120] = 8'hce ;
            rom[13121] = 8'h04 ;
            rom[13122] = 8'hf4 ;
            rom[13123] = 8'h20 ;
            rom[13124] = 8'h0f ;
            rom[13125] = 8'h3c ;
            rom[13126] = 8'hb7 ;
            rom[13127] = 8'h05 ;
            rom[13128] = 8'h1d ;
            rom[13129] = 8'hf9 ;
            rom[13130] = 8'h08 ;
            rom[13131] = 8'h04 ;
            rom[13132] = 8'h10 ;
            rom[13133] = 8'hc6 ;
            rom[13134] = 8'h26 ;
            rom[13135] = 8'hfd ;
            rom[13136] = 8'hf2 ;
            rom[13137] = 8'h01 ;
            rom[13138] = 8'h05 ;
            rom[13139] = 8'hf2 ;
            rom[13140] = 8'he7 ;
            rom[13141] = 8'h12 ;
            rom[13142] = 8'hf5 ;
            rom[13143] = 8'hea ;
            rom[13144] = 8'hff ;
            rom[13145] = 8'hde ;
            rom[13146] = 8'hfd ;
            rom[13147] = 8'hfa ;
            rom[13148] = 8'h2b ;
            rom[13149] = 8'he9 ;
            rom[13150] = 8'h0d ;
            rom[13151] = 8'h00 ;
            rom[13152] = 8'h12 ;
            rom[13153] = 8'hfa ;
            rom[13154] = 8'hfb ;
            rom[13155] = 8'h0b ;
            rom[13156] = 8'h24 ;
            rom[13157] = 8'hfc ;
            rom[13158] = 8'h15 ;
            rom[13159] = 8'hfd ;
            rom[13160] = 8'hf7 ;
            rom[13161] = 8'h0a ;
            rom[13162] = 8'hfb ;
            rom[13163] = 8'h17 ;
            rom[13164] = 8'h13 ;
            rom[13165] = 8'h16 ;
            rom[13166] = 8'he4 ;
            rom[13167] = 8'he5 ;
            rom[13168] = 8'hec ;
            rom[13169] = 8'h03 ;
            rom[13170] = 8'h07 ;
            rom[13171] = 8'h12 ;
            rom[13172] = 8'h0d ;
            rom[13173] = 8'h11 ;
            rom[13174] = 8'hf3 ;
            rom[13175] = 8'hf2 ;
            rom[13176] = 8'hf1 ;
            rom[13177] = 8'hd9 ;
            rom[13178] = 8'h10 ;
            rom[13179] = 8'hf6 ;
            rom[13180] = 8'h02 ;
            rom[13181] = 8'h25 ;
            rom[13182] = 8'h1f ;
            rom[13183] = 8'h0e ;
            rom[13184] = 8'h0e ;
            rom[13185] = 8'hfb ;
            rom[13186] = 8'h23 ;
            rom[13187] = 8'hdd ;
            rom[13188] = 8'hff ;
            rom[13189] = 8'h0e ;
            rom[13190] = 8'he4 ;
            rom[13191] = 8'hfc ;
            rom[13192] = 8'h32 ;
            rom[13193] = 8'hf5 ;
            rom[13194] = 8'hf1 ;
            rom[13195] = 8'h20 ;
            rom[13196] = 8'h0b ;
            rom[13197] = 8'hde ;
            rom[13198] = 8'hfe ;
            rom[13199] = 8'h13 ;
            rom[13200] = 8'h10 ;
            rom[13201] = 8'h1d ;
            rom[13202] = 8'h04 ;
            rom[13203] = 8'h16 ;
            rom[13204] = 8'h07 ;
            rom[13205] = 8'hf4 ;
            rom[13206] = 8'hf7 ;
            rom[13207] = 8'hfd ;
            rom[13208] = 8'hdc ;
            rom[13209] = 8'hfb ;
            rom[13210] = 8'h20 ;
            rom[13211] = 8'hfb ;
            rom[13212] = 8'hda ;
            rom[13213] = 8'h0c ;
            rom[13214] = 8'hf8 ;
            rom[13215] = 8'he4 ;
            rom[13216] = 8'hee ;
            rom[13217] = 8'h14 ;
            rom[13218] = 8'hfe ;
            rom[13219] = 8'hda ;
            rom[13220] = 8'hed ;
            rom[13221] = 8'hf9 ;
            rom[13222] = 8'h16 ;
            rom[13223] = 8'hbd ;
            rom[13224] = 8'hf9 ;
            rom[13225] = 8'hf5 ;
            rom[13226] = 8'hff ;
            rom[13227] = 8'h25 ;
            rom[13228] = 8'h0a ;
            rom[13229] = 8'hf7 ;
            rom[13230] = 8'h00 ;
            rom[13231] = 8'h0e ;
            rom[13232] = 8'hed ;
            rom[13233] = 8'he6 ;
            rom[13234] = 8'h03 ;
            rom[13235] = 8'hfe ;
            rom[13236] = 8'hfe ;
            rom[13237] = 8'hdb ;
            rom[13238] = 8'hf7 ;
            rom[13239] = 8'h01 ;
            rom[13240] = 8'hfd ;
            rom[13241] = 8'he7 ;
            rom[13242] = 8'h27 ;
            rom[13243] = 8'hc9 ;
            rom[13244] = 8'he7 ;
            rom[13245] = 8'hdc ;
            rom[13246] = 8'h13 ;
            rom[13247] = 8'hf7 ;
            rom[13248] = 8'he8 ;
            rom[13249] = 8'hf6 ;
            rom[13250] = 8'hed ;
            rom[13251] = 8'hfb ;
            rom[13252] = 8'hf9 ;
            rom[13253] = 8'hfa ;
            rom[13254] = 8'hfd ;
            rom[13255] = 8'h07 ;
            rom[13256] = 8'hfa ;
            rom[13257] = 8'hfe ;
            rom[13258] = 8'h14 ;
            rom[13259] = 8'h06 ;
            rom[13260] = 8'hff ;
            rom[13261] = 8'h02 ;
            rom[13262] = 8'h14 ;
            rom[13263] = 8'hd7 ;
            rom[13264] = 8'hed ;
            rom[13265] = 8'h05 ;
            rom[13266] = 8'hf0 ;
            rom[13267] = 8'he5 ;
            rom[13268] = 8'h18 ;
            rom[13269] = 8'hd3 ;
            rom[13270] = 8'hf2 ;
            rom[13271] = 8'h2c ;
            rom[13272] = 8'h02 ;
            rom[13273] = 8'hf3 ;
            rom[13274] = 8'h0f ;
            rom[13275] = 8'hfc ;
            rom[13276] = 8'h10 ;
            rom[13277] = 8'he5 ;
            rom[13278] = 8'h00 ;
            rom[13279] = 8'hf5 ;
            rom[13280] = 8'h06 ;
            rom[13281] = 8'h22 ;
            rom[13282] = 8'he2 ;
            rom[13283] = 8'h02 ;
            rom[13284] = 8'he8 ;
            rom[13285] = 8'hde ;
            rom[13286] = 8'hf0 ;
            rom[13287] = 8'hfe ;
            rom[13288] = 8'h0c ;
            rom[13289] = 8'h1a ;
            rom[13290] = 8'h09 ;
            rom[13291] = 8'h01 ;
            rom[13292] = 8'h00 ;
            rom[13293] = 8'h0e ;
            rom[13294] = 8'hf0 ;
            rom[13295] = 8'hd8 ;
            rom[13296] = 8'hce ;
            rom[13297] = 8'hed ;
            rom[13298] = 8'heb ;
            rom[13299] = 8'h09 ;
            rom[13300] = 8'hfb ;
            rom[13301] = 8'h00 ;
            rom[13302] = 8'h11 ;
            rom[13303] = 8'h36 ;
            rom[13304] = 8'h0b ;
            rom[13305] = 8'h09 ;
            rom[13306] = 8'he1 ;
            rom[13307] = 8'hd8 ;
            rom[13308] = 8'h23 ;
            rom[13309] = 8'hfa ;
            rom[13310] = 8'h15 ;
            rom[13311] = 8'he3 ;
            rom[13312] = 8'h21 ;
            rom[13313] = 8'hf7 ;
            rom[13314] = 8'h10 ;
            rom[13315] = 8'h1a ;
            rom[13316] = 8'hf2 ;
            rom[13317] = 8'hb0 ;
            rom[13318] = 8'h04 ;
            rom[13319] = 8'h14 ;
            rom[13320] = 8'h1e ;
            rom[13321] = 8'he1 ;
            rom[13322] = 8'hec ;
            rom[13323] = 8'hff ;
            rom[13324] = 8'hee ;
            rom[13325] = 8'hfb ;
            rom[13326] = 8'hf1 ;
            rom[13327] = 8'hdb ;
            rom[13328] = 8'hf6 ;
            rom[13329] = 8'hd9 ;
            rom[13330] = 8'h11 ;
            rom[13331] = 8'h0b ;
            rom[13332] = 8'h00 ;
            rom[13333] = 8'he8 ;
            rom[13334] = 8'hed ;
            rom[13335] = 8'hca ;
            rom[13336] = 8'hf8 ;
            rom[13337] = 8'h04 ;
            rom[13338] = 8'hdd ;
            rom[13339] = 8'h09 ;
            rom[13340] = 8'h01 ;
            rom[13341] = 8'h10 ;
            rom[13342] = 8'h16 ;
            rom[13343] = 8'he8 ;
            rom[13344] = 8'hdf ;
            rom[13345] = 8'hfa ;
            rom[13346] = 8'h0a ;
            rom[13347] = 8'hdf ;
            rom[13348] = 8'hf4 ;
            rom[13349] = 8'h05 ;
            rom[13350] = 8'h02 ;
            rom[13351] = 8'hf8 ;
            rom[13352] = 8'hee ;
            rom[13353] = 8'hf5 ;
            rom[13354] = 8'hfa ;
            rom[13355] = 8'hf4 ;
            rom[13356] = 8'h0e ;
            rom[13357] = 8'h09 ;
            rom[13358] = 8'hd0 ;
            rom[13359] = 8'h1f ;
            rom[13360] = 8'h02 ;
            rom[13361] = 8'h07 ;
            rom[13362] = 8'hfc ;
            rom[13363] = 8'hf5 ;
            rom[13364] = 8'h14 ;
            rom[13365] = 8'hf4 ;
            rom[13366] = 8'heb ;
            rom[13367] = 8'h00 ;
            rom[13368] = 8'h0e ;
            rom[13369] = 8'hf3 ;
            rom[13370] = 8'hf2 ;
            rom[13371] = 8'hd9 ;
            rom[13372] = 8'hf1 ;
            rom[13373] = 8'h0a ;
            rom[13374] = 8'hd9 ;
            rom[13375] = 8'h1c ;
            rom[13376] = 8'h0d ;
            rom[13377] = 8'h0f ;
            rom[13378] = 8'hee ;
            rom[13379] = 8'hd5 ;
            rom[13380] = 8'h06 ;
            rom[13381] = 8'h00 ;
            rom[13382] = 8'h02 ;
            rom[13383] = 8'hd7 ;
            rom[13384] = 8'he4 ;
            rom[13385] = 8'hf2 ;
            rom[13386] = 8'hf9 ;
            rom[13387] = 8'h0a ;
            rom[13388] = 8'h04 ;
            rom[13389] = 8'h06 ;
            rom[13390] = 8'hdb ;
            rom[13391] = 8'hf7 ;
            rom[13392] = 8'h06 ;
            rom[13393] = 8'hf7 ;
            rom[13394] = 8'hee ;
            rom[13395] = 8'h1a ;
            rom[13396] = 8'hf2 ;
            rom[13397] = 8'h12 ;
            rom[13398] = 8'h03 ;
            rom[13399] = 8'hf7 ;
            rom[13400] = 8'hf3 ;
            rom[13401] = 8'hd3 ;
            rom[13402] = 8'hfb ;
            rom[13403] = 8'he5 ;
            rom[13404] = 8'hcf ;
            rom[13405] = 8'h04 ;
            rom[13406] = 8'hf7 ;
            rom[13407] = 8'he0 ;
            rom[13408] = 8'hf3 ;
            rom[13409] = 8'hff ;
            rom[13410] = 8'hf0 ;
            rom[13411] = 8'h19 ;
            rom[13412] = 8'hfc ;
            rom[13413] = 8'h03 ;
            rom[13414] = 8'hff ;
            rom[13415] = 8'hfa ;
            rom[13416] = 8'hc4 ;
            rom[13417] = 8'hdc ;
            rom[13418] = 8'hec ;
            rom[13419] = 8'hf5 ;
            rom[13420] = 8'hec ;
            rom[13421] = 8'h2a ;
            rom[13422] = 8'h03 ;
            rom[13423] = 8'h2c ;
            rom[13424] = 8'h04 ;
            rom[13425] = 8'hd9 ;
            rom[13426] = 8'h16 ;
            rom[13427] = 8'h07 ;
            rom[13428] = 8'hdc ;
            rom[13429] = 8'hd2 ;
            rom[13430] = 8'hca ;
            rom[13431] = 8'hc9 ;
            rom[13432] = 8'hf5 ;
            rom[13433] = 8'he2 ;
            rom[13434] = 8'hef ;
            rom[13435] = 8'h03 ;
            rom[13436] = 8'hea ;
            rom[13437] = 8'hc7 ;
            rom[13438] = 8'hf1 ;
            rom[13439] = 8'h17 ;
            rom[13440] = 8'h08 ;
            rom[13441] = 8'hf8 ;
            rom[13442] = 8'h10 ;
            rom[13443] = 8'h10 ;
            rom[13444] = 8'hfa ;
            rom[13445] = 8'h01 ;
            rom[13446] = 8'hf9 ;
            rom[13447] = 8'he1 ;
            rom[13448] = 8'hee ;
            rom[13449] = 8'h0a ;
            rom[13450] = 8'hdd ;
            rom[13451] = 8'h03 ;
            rom[13452] = 8'he5 ;
            rom[13453] = 8'h07 ;
            rom[13454] = 8'hf4 ;
            rom[13455] = 8'h0f ;
            rom[13456] = 8'hf4 ;
            rom[13457] = 8'h1f ;
            rom[13458] = 8'hd7 ;
            rom[13459] = 8'h02 ;
            rom[13460] = 8'h0a ;
            rom[13461] = 8'h06 ;
            rom[13462] = 8'hb5 ;
            rom[13463] = 8'hf6 ;
            rom[13464] = 8'hec ;
            rom[13465] = 8'h04 ;
            rom[13466] = 8'h0f ;
            rom[13467] = 8'hf0 ;
            rom[13468] = 8'hf5 ;
            rom[13469] = 8'h0a ;
            rom[13470] = 8'h09 ;
            rom[13471] = 8'h0d ;
            rom[13472] = 8'he9 ;
            rom[13473] = 8'h1a ;
            rom[13474] = 8'h07 ;
            rom[13475] = 8'h09 ;
            rom[13476] = 8'hf6 ;
            rom[13477] = 8'he9 ;
            rom[13478] = 8'hfa ;
            rom[13479] = 8'hfa ;
            rom[13480] = 8'hf0 ;
            rom[13481] = 8'he8 ;
            rom[13482] = 8'hf2 ;
            rom[13483] = 8'hf3 ;
            rom[13484] = 8'hf0 ;
            rom[13485] = 8'he4 ;
            rom[13486] = 8'hf4 ;
            rom[13487] = 8'hf6 ;
            rom[13488] = 8'hb7 ;
            rom[13489] = 8'hc4 ;
            rom[13490] = 8'hf6 ;
            rom[13491] = 8'hed ;
            rom[13492] = 8'hf9 ;
            rom[13493] = 8'hf8 ;
            rom[13494] = 8'hc6 ;
            rom[13495] = 8'h15 ;
            rom[13496] = 8'h06 ;
            rom[13497] = 8'hef ;
            rom[13498] = 8'h07 ;
            rom[13499] = 8'hc0 ;
            rom[13500] = 8'he0 ;
            rom[13501] = 8'hc2 ;
            rom[13502] = 8'h1c ;
            rom[13503] = 8'hfd ;
            rom[13504] = 8'hcd ;
            rom[13505] = 8'h0e ;
            rom[13506] = 8'hd9 ;
            rom[13507] = 8'h3c ;
            rom[13508] = 8'hf2 ;
            rom[13509] = 8'he0 ;
            rom[13510] = 8'hf7 ;
            rom[13511] = 8'h06 ;
            rom[13512] = 8'hf3 ;
            rom[13513] = 8'h0c ;
            rom[13514] = 8'h0a ;
            rom[13515] = 8'h10 ;
            rom[13516] = 8'h03 ;
            rom[13517] = 8'h04 ;
            rom[13518] = 8'h27 ;
            rom[13519] = 8'h0b ;
            rom[13520] = 8'hd2 ;
            rom[13521] = 8'hff ;
            rom[13522] = 8'hd2 ;
            rom[13523] = 8'h13 ;
            rom[13524] = 8'he8 ;
            rom[13525] = 8'hf6 ;
            rom[13526] = 8'hf1 ;
            rom[13527] = 8'hfd ;
            rom[13528] = 8'h04 ;
            rom[13529] = 8'h02 ;
            rom[13530] = 8'h0a ;
            rom[13531] = 8'h0d ;
            rom[13532] = 8'h30 ;
            rom[13533] = 8'h14 ;
            rom[13534] = 8'h0c ;
            rom[13535] = 8'h07 ;
            rom[13536] = 8'hfa ;
            rom[13537] = 8'hd5 ;
            rom[13538] = 8'h22 ;
            rom[13539] = 8'hc4 ;
            rom[13540] = 8'hdf ;
            rom[13541] = 8'hf1 ;
            rom[13542] = 8'he9 ;
            rom[13543] = 8'h06 ;
            rom[13544] = 8'hfb ;
            rom[13545] = 8'hef ;
            rom[13546] = 8'hf3 ;
            rom[13547] = 8'hf3 ;
            rom[13548] = 8'hfa ;
            rom[13549] = 8'h07 ;
            rom[13550] = 8'hf4 ;
            rom[13551] = 8'h02 ;
            rom[13552] = 8'he6 ;
            rom[13553] = 8'he9 ;
            rom[13554] = 8'h1c ;
            rom[13555] = 8'h31 ;
            rom[13556] = 8'h09 ;
            rom[13557] = 8'hf6 ;
            rom[13558] = 8'hfd ;
            rom[13559] = 8'h03 ;
            rom[13560] = 8'he1 ;
            rom[13561] = 8'hef ;
            rom[13562] = 8'hf5 ;
            rom[13563] = 8'he9 ;
            rom[13564] = 8'h13 ;
            rom[13565] = 8'hfe ;
            rom[13566] = 8'hfe ;
            rom[13567] = 8'h03 ;
            rom[13568] = 8'hdd ;
            rom[13569] = 8'h02 ;
            rom[13570] = 8'he6 ;
            rom[13571] = 8'he4 ;
            rom[13572] = 8'h06 ;
            rom[13573] = 8'h08 ;
            rom[13574] = 8'he6 ;
            rom[13575] = 8'h0c ;
            rom[13576] = 8'h0d ;
            rom[13577] = 8'hcc ;
            rom[13578] = 8'hfa ;
            rom[13579] = 8'he6 ;
            rom[13580] = 8'hf6 ;
            rom[13581] = 8'hf7 ;
            rom[13582] = 8'h04 ;
            rom[13583] = 8'hdb ;
            rom[13584] = 8'h0c ;
            rom[13585] = 8'he6 ;
            rom[13586] = 8'hd8 ;
            rom[13587] = 8'hff ;
            rom[13588] = 8'hfe ;
            rom[13589] = 8'h02 ;
            rom[13590] = 8'h12 ;
            rom[13591] = 8'hff ;
            rom[13592] = 8'h0d ;
            rom[13593] = 8'hf7 ;
            rom[13594] = 8'h1e ;
            rom[13595] = 8'h04 ;
            rom[13596] = 8'h24 ;
            rom[13597] = 8'h03 ;
            rom[13598] = 8'hec ;
            rom[13599] = 8'hdf ;
            rom[13600] = 8'h32 ;
            rom[13601] = 8'hef ;
            rom[13602] = 8'hd7 ;
            rom[13603] = 8'h00 ;
            rom[13604] = 8'hed ;
            rom[13605] = 8'h01 ;
            rom[13606] = 8'h17 ;
            rom[13607] = 8'h0f ;
            rom[13608] = 8'hf3 ;
            rom[13609] = 8'hce ;
            rom[13610] = 8'hf1 ;
            rom[13611] = 8'h02 ;
            rom[13612] = 8'h24 ;
            rom[13613] = 8'h23 ;
            rom[13614] = 8'h00 ;
            rom[13615] = 8'he7 ;
            rom[13616] = 8'hea ;
            rom[13617] = 8'h0f ;
            rom[13618] = 8'h05 ;
            rom[13619] = 8'hfe ;
            rom[13620] = 8'hf2 ;
            rom[13621] = 8'h02 ;
            rom[13622] = 8'h0e ;
            rom[13623] = 8'h04 ;
            rom[13624] = 8'hf3 ;
            rom[13625] = 8'hec ;
            rom[13626] = 8'h0a ;
            rom[13627] = 8'hc7 ;
            rom[13628] = 8'he3 ;
            rom[13629] = 8'hfd ;
            rom[13630] = 8'he7 ;
            rom[13631] = 8'h0d ;
            rom[13632] = 8'h01 ;
            rom[13633] = 8'hba ;
            rom[13634] = 8'h00 ;
            rom[13635] = 8'h0d ;
            rom[13636] = 8'hf5 ;
            rom[13637] = 8'hf3 ;
            rom[13638] = 8'h24 ;
            rom[13639] = 8'hf5 ;
            rom[13640] = 8'he9 ;
            rom[13641] = 8'hc3 ;
            rom[13642] = 8'hfb ;
            rom[13643] = 8'h00 ;
            rom[13644] = 8'h07 ;
            rom[13645] = 8'hcf ;
            rom[13646] = 8'hc8 ;
            rom[13647] = 8'h08 ;
            rom[13648] = 8'h1d ;
            rom[13649] = 8'hdf ;
            rom[13650] = 8'h1a ;
            rom[13651] = 8'he7 ;
            rom[13652] = 8'hed ;
            rom[13653] = 8'h05 ;
            rom[13654] = 8'hee ;
            rom[13655] = 8'hdf ;
            rom[13656] = 8'hf8 ;
            rom[13657] = 8'hfd ;
            rom[13658] = 8'h02 ;
            rom[13659] = 8'h13 ;
            rom[13660] = 8'h13 ;
            rom[13661] = 8'h0d ;
            rom[13662] = 8'h08 ;
            rom[13663] = 8'hf0 ;
            rom[13664] = 8'hfd ;
            rom[13665] = 8'h04 ;
            rom[13666] = 8'hfb ;
            rom[13667] = 8'he4 ;
            rom[13668] = 8'h0a ;
            rom[13669] = 8'hef ;
            rom[13670] = 8'h0d ;
            rom[13671] = 8'hfd ;
            rom[13672] = 8'hfd ;
            rom[13673] = 8'hed ;
            rom[13674] = 8'h20 ;
            rom[13675] = 8'h18 ;
            rom[13676] = 8'h01 ;
            rom[13677] = 8'h12 ;
            rom[13678] = 8'hdf ;
            rom[13679] = 8'he4 ;
            rom[13680] = 8'h0e ;
            rom[13681] = 8'hf7 ;
            rom[13682] = 8'h2a ;
            rom[13683] = 8'h00 ;
            rom[13684] = 8'hf2 ;
            rom[13685] = 8'he4 ;
            rom[13686] = 8'h02 ;
            rom[13687] = 8'h0b ;
            rom[13688] = 8'hd3 ;
            rom[13689] = 8'hf2 ;
            rom[13690] = 8'h14 ;
            rom[13691] = 8'hf5 ;
            rom[13692] = 8'h08 ;
            rom[13693] = 8'h0b ;
            rom[13694] = 8'h12 ;
            rom[13695] = 8'hfc ;
            rom[13696] = 8'he1 ;
            rom[13697] = 8'h11 ;
            rom[13698] = 8'hf2 ;
            rom[13699] = 8'h0f ;
            rom[13700] = 8'hf8 ;
            rom[13701] = 8'hdd ;
            rom[13702] = 8'hfc ;
            rom[13703] = 8'h04 ;
            rom[13704] = 8'hfd ;
            rom[13705] = 8'hdf ;
            rom[13706] = 8'h18 ;
            rom[13707] = 8'hee ;
            rom[13708] = 8'hfb ;
            rom[13709] = 8'hf1 ;
            rom[13710] = 8'hd9 ;
            rom[13711] = 8'h01 ;
            rom[13712] = 8'he4 ;
            rom[13713] = 8'hd4 ;
            rom[13714] = 8'hf8 ;
            rom[13715] = 8'hde ;
            rom[13716] = 8'h1a ;
            rom[13717] = 8'h27 ;
            rom[13718] = 8'h00 ;
            rom[13719] = 8'hfc ;
            rom[13720] = 8'he5 ;
            rom[13721] = 8'he8 ;
            rom[13722] = 8'heb ;
            rom[13723] = 8'hfe ;
            rom[13724] = 8'hfc ;
            rom[13725] = 8'hf1 ;
            rom[13726] = 8'h0f ;
            rom[13727] = 8'he0 ;
            rom[13728] = 8'hfc ;
            rom[13729] = 8'h13 ;
            rom[13730] = 8'hcd ;
            rom[13731] = 8'h03 ;
            rom[13732] = 8'hfa ;
            rom[13733] = 8'hfd ;
            rom[13734] = 8'h00 ;
            rom[13735] = 8'h00 ;
            rom[13736] = 8'hf8 ;
            rom[13737] = 8'hea ;
            rom[13738] = 8'h16 ;
            rom[13739] = 8'hf7 ;
            rom[13740] = 8'hf5 ;
            rom[13741] = 8'hf6 ;
            rom[13742] = 8'h11 ;
            rom[13743] = 8'h1e ;
            rom[13744] = 8'hff ;
            rom[13745] = 8'hf0 ;
            rom[13746] = 8'hed ;
            rom[13747] = 8'h12 ;
            rom[13748] = 8'h0f ;
            rom[13749] = 8'h10 ;
            rom[13750] = 8'he6 ;
            rom[13751] = 8'h27 ;
            rom[13752] = 8'hfb ;
            rom[13753] = 8'h04 ;
            rom[13754] = 8'he7 ;
            rom[13755] = 8'hfd ;
            rom[13756] = 8'hfc ;
            rom[13757] = 8'h06 ;
            rom[13758] = 8'hc2 ;
            rom[13759] = 8'he2 ;
            rom[13760] = 8'h04 ;
            rom[13761] = 8'he1 ;
            rom[13762] = 8'hf4 ;
            rom[13763] = 8'h19 ;
            rom[13764] = 8'he8 ;
            rom[13765] = 8'hf9 ;
            rom[13766] = 8'h15 ;
            rom[13767] = 8'h03 ;
            rom[13768] = 8'hf7 ;
            rom[13769] = 8'hc9 ;
            rom[13770] = 8'h13 ;
            rom[13771] = 8'hfe ;
            rom[13772] = 8'hfb ;
            rom[13773] = 8'h01 ;
            rom[13774] = 8'hd0 ;
            rom[13775] = 8'he7 ;
            rom[13776] = 8'h01 ;
            rom[13777] = 8'heb ;
            rom[13778] = 8'hd4 ;
            rom[13779] = 8'h16 ;
            rom[13780] = 8'hde ;
            rom[13781] = 8'hd8 ;
            rom[13782] = 8'hf6 ;
            rom[13783] = 8'h14 ;
            rom[13784] = 8'h06 ;
            rom[13785] = 8'h08 ;
            rom[13786] = 8'h0c ;
            rom[13787] = 8'h05 ;
            rom[13788] = 8'hea ;
            rom[13789] = 8'he5 ;
            rom[13790] = 8'heb ;
            rom[13791] = 8'hfd ;
            rom[13792] = 8'heb ;
            rom[13793] = 8'h23 ;
            rom[13794] = 8'hd5 ;
            rom[13795] = 8'hfc ;
            rom[13796] = 8'hf7 ;
            rom[13797] = 8'hfd ;
            rom[13798] = 8'hf1 ;
            rom[13799] = 8'he9 ;
            rom[13800] = 8'hfa ;
            rom[13801] = 8'hdc ;
            rom[13802] = 8'he9 ;
            rom[13803] = 8'hf5 ;
            rom[13804] = 8'he1 ;
            rom[13805] = 8'h01 ;
            rom[13806] = 8'hd1 ;
            rom[13807] = 8'h2a ;
            rom[13808] = 8'hee ;
            rom[13809] = 8'he7 ;
            rom[13810] = 8'h19 ;
            rom[13811] = 8'h10 ;
            rom[13812] = 8'hea ;
            rom[13813] = 8'h00 ;
            rom[13814] = 8'hef ;
            rom[13815] = 8'hca ;
            rom[13816] = 8'hfd ;
            rom[13817] = 8'h0d ;
            rom[13818] = 8'hf3 ;
            rom[13819] = 8'hf2 ;
            rom[13820] = 8'h22 ;
            rom[13821] = 8'hdc ;
            rom[13822] = 8'hf5 ;
            rom[13823] = 8'hf8 ;
            rom[13824] = 8'hf6 ;
            rom[13825] = 8'hcd ;
            rom[13826] = 8'h18 ;
            rom[13827] = 8'hf7 ;
            rom[13828] = 8'he3 ;
            rom[13829] = 8'hf9 ;
            rom[13830] = 8'hdc ;
            rom[13831] = 8'he2 ;
            rom[13832] = 8'hef ;
            rom[13833] = 8'hc5 ;
            rom[13834] = 8'hf6 ;
            rom[13835] = 8'h1b ;
            rom[13836] = 8'hfb ;
            rom[13837] = 8'h09 ;
            rom[13838] = 8'h0d ;
            rom[13839] = 8'hd4 ;
            rom[13840] = 8'he4 ;
            rom[13841] = 8'h18 ;
            rom[13842] = 8'hda ;
            rom[13843] = 8'h20 ;
            rom[13844] = 8'hf9 ;
            rom[13845] = 8'he2 ;
            rom[13846] = 8'h31 ;
            rom[13847] = 8'hec ;
            rom[13848] = 8'hf4 ;
            rom[13849] = 8'hbc ;
            rom[13850] = 8'h0c ;
            rom[13851] = 8'haf ;
            rom[13852] = 8'hec ;
            rom[13853] = 8'hcf ;
            rom[13854] = 8'hf1 ;
            rom[13855] = 8'hea ;
            rom[13856] = 8'h14 ;
            rom[13857] = 8'h25 ;
            rom[13858] = 8'h05 ;
            rom[13859] = 8'he6 ;
            rom[13860] = 8'h06 ;
            rom[13861] = 8'h02 ;
            rom[13862] = 8'h0b ;
            rom[13863] = 8'he0 ;
            rom[13864] = 8'h1e ;
            rom[13865] = 8'hda ;
            rom[13866] = 8'hf8 ;
            rom[13867] = 8'he3 ;
            rom[13868] = 8'hcf ;
            rom[13869] = 8'he7 ;
            rom[13870] = 8'hf2 ;
            rom[13871] = 8'h05 ;
            rom[13872] = 8'h01 ;
            rom[13873] = 8'hda ;
            rom[13874] = 8'hfd ;
            rom[13875] = 8'hfd ;
            rom[13876] = 8'hfe ;
            rom[13877] = 8'h09 ;
            rom[13878] = 8'h00 ;
            rom[13879] = 8'hfb ;
            rom[13880] = 8'hf5 ;
            rom[13881] = 8'hda ;
            rom[13882] = 8'hd9 ;
            rom[13883] = 8'he3 ;
            rom[13884] = 8'he4 ;
            rom[13885] = 8'hf0 ;
            rom[13886] = 8'h03 ;
            rom[13887] = 8'hcd ;
            rom[13888] = 8'hce ;
            rom[13889] = 8'hed ;
            rom[13890] = 8'h04 ;
            rom[13891] = 8'hfc ;
            rom[13892] = 8'h0d ;
            rom[13893] = 8'h09 ;
            rom[13894] = 8'hee ;
            rom[13895] = 8'h21 ;
            rom[13896] = 8'h06 ;
            rom[13897] = 8'hfc ;
            rom[13898] = 8'hf3 ;
            rom[13899] = 8'heb ;
            rom[13900] = 8'hc7 ;
            rom[13901] = 8'h07 ;
            rom[13902] = 8'hf4 ;
            rom[13903] = 8'he4 ;
            rom[13904] = 8'he9 ;
            rom[13905] = 8'heb ;
            rom[13906] = 8'h1c ;
            rom[13907] = 8'hd9 ;
            rom[13908] = 8'h00 ;
            rom[13909] = 8'hd9 ;
            rom[13910] = 8'h00 ;
            rom[13911] = 8'hfa ;
            rom[13912] = 8'hd8 ;
            rom[13913] = 8'hf8 ;
            rom[13914] = 8'h0c ;
            rom[13915] = 8'h16 ;
            rom[13916] = 8'hee ;
            rom[13917] = 8'hdc ;
            rom[13918] = 8'h12 ;
            rom[13919] = 8'hff ;
            rom[13920] = 8'h0b ;
            rom[13921] = 8'h03 ;
            rom[13922] = 8'hfa ;
            rom[13923] = 8'h18 ;
            rom[13924] = 8'he0 ;
            rom[13925] = 8'hf5 ;
            rom[13926] = 8'he5 ;
            rom[13927] = 8'hed ;
            rom[13928] = 8'he9 ;
            rom[13929] = 8'h16 ;
            rom[13930] = 8'he0 ;
            rom[13931] = 8'hf1 ;
            rom[13932] = 8'hfa ;
            rom[13933] = 8'h0b ;
            rom[13934] = 8'hf3 ;
            rom[13935] = 8'h22 ;
            rom[13936] = 8'hf3 ;
            rom[13937] = 8'h22 ;
            rom[13938] = 8'h07 ;
            rom[13939] = 8'he9 ;
            rom[13940] = 8'hd1 ;
            rom[13941] = 8'h04 ;
            rom[13942] = 8'hfd ;
            rom[13943] = 8'h14 ;
            rom[13944] = 8'h04 ;
            rom[13945] = 8'h00 ;
            rom[13946] = 8'hf0 ;
            rom[13947] = 8'hee ;
            rom[13948] = 8'hf1 ;
            rom[13949] = 8'hfe ;
            rom[13950] = 8'he2 ;
            rom[13951] = 8'h1a ;
            rom[13952] = 8'h03 ;
            rom[13953] = 8'hef ;
            rom[13954] = 8'h05 ;
            rom[13955] = 8'h0b ;
            rom[13956] = 8'hf9 ;
            rom[13957] = 8'hbe ;
            rom[13958] = 8'hf2 ;
            rom[13959] = 8'h14 ;
            rom[13960] = 8'hec ;
            rom[13961] = 8'hdc ;
            rom[13962] = 8'h04 ;
            rom[13963] = 8'h0d ;
            rom[13964] = 8'hf1 ;
            rom[13965] = 8'he6 ;
            rom[13966] = 8'h0b ;
            rom[13967] = 8'h0f ;
            rom[13968] = 8'hef ;
            rom[13969] = 8'hdd ;
            rom[13970] = 8'he4 ;
            rom[13971] = 8'hdb ;
            rom[13972] = 8'h03 ;
            rom[13973] = 8'he6 ;
            rom[13974] = 8'h07 ;
            rom[13975] = 8'hf9 ;
            rom[13976] = 8'he3 ;
            rom[13977] = 8'hda ;
            rom[13978] = 8'h06 ;
            rom[13979] = 8'he1 ;
            rom[13980] = 8'h00 ;
            rom[13981] = 8'hd9 ;
            rom[13982] = 8'h05 ;
            rom[13983] = 8'hf2 ;
            rom[13984] = 8'h0c ;
            rom[13985] = 8'h10 ;
            rom[13986] = 8'h03 ;
            rom[13987] = 8'hcc ;
            rom[13988] = 8'he3 ;
            rom[13989] = 8'hfd ;
            rom[13990] = 8'h11 ;
            rom[13991] = 8'h00 ;
            rom[13992] = 8'hd3 ;
            rom[13993] = 8'h05 ;
            rom[13994] = 8'h35 ;
            rom[13995] = 8'hcf ;
            rom[13996] = 8'hdc ;
            rom[13997] = 8'h21 ;
            rom[13998] = 8'hd0 ;
            rom[13999] = 8'hfe ;
            rom[14000] = 8'h1e ;
            rom[14001] = 8'hdd ;
            rom[14002] = 8'hff ;
            rom[14003] = 8'hf0 ;
            rom[14004] = 8'h12 ;
            rom[14005] = 8'h0c ;
            rom[14006] = 8'hdf ;
            rom[14007] = 8'hf7 ;
            rom[14008] = 8'hde ;
            rom[14009] = 8'hef ;
            rom[14010] = 8'hdf ;
            rom[14011] = 8'h15 ;
            rom[14012] = 8'h0a ;
            rom[14013] = 8'h10 ;
            rom[14014] = 8'hda ;
            rom[14015] = 8'hd1 ;
            rom[14016] = 8'hef ;
            rom[14017] = 8'hfd ;
            rom[14018] = 8'hfb ;
            rom[14019] = 8'hfd ;
            rom[14020] = 8'hfb ;
            rom[14021] = 8'hfe ;
            rom[14022] = 8'h04 ;
            rom[14023] = 8'h0f ;
            rom[14024] = 8'h21 ;
            rom[14025] = 8'hd3 ;
            rom[14026] = 8'he1 ;
            rom[14027] = 8'he5 ;
            rom[14028] = 8'h0f ;
            rom[14029] = 8'hf4 ;
            rom[14030] = 8'hf3 ;
            rom[14031] = 8'hed ;
            rom[14032] = 8'hf2 ;
            rom[14033] = 8'he6 ;
            rom[14034] = 8'he8 ;
            rom[14035] = 8'h00 ;
            rom[14036] = 8'hfd ;
            rom[14037] = 8'hdf ;
            rom[14038] = 8'h01 ;
            rom[14039] = 8'h0a ;
            rom[14040] = 8'h08 ;
            rom[14041] = 8'h0d ;
            rom[14042] = 8'h0e ;
            rom[14043] = 8'h0c ;
            rom[14044] = 8'hd1 ;
            rom[14045] = 8'hd4 ;
            rom[14046] = 8'h0d ;
            rom[14047] = 8'hf6 ;
            rom[14048] = 8'hdc ;
            rom[14049] = 8'h0d ;
            rom[14050] = 8'hcf ;
            rom[14051] = 8'hfd ;
            rom[14052] = 8'hdf ;
            rom[14053] = 8'h21 ;
            rom[14054] = 8'h11 ;
            rom[14055] = 8'hf0 ;
            rom[14056] = 8'hf6 ;
            rom[14057] = 8'h00 ;
            rom[14058] = 8'h05 ;
            rom[14059] = 8'he1 ;
            rom[14060] = 8'hff ;
            rom[14061] = 8'h0a ;
            rom[14062] = 8'h04 ;
            rom[14063] = 8'h20 ;
            rom[14064] = 8'he3 ;
            rom[14065] = 8'h0c ;
            rom[14066] = 8'h10 ;
            rom[14067] = 8'hf5 ;
            rom[14068] = 8'hcd ;
            rom[14069] = 8'h06 ;
            rom[14070] = 8'hf1 ;
            rom[14071] = 8'h0c ;
            rom[14072] = 8'h03 ;
            rom[14073] = 8'he9 ;
            rom[14074] = 8'hed ;
            rom[14075] = 8'hf2 ;
            rom[14076] = 8'hf1 ;
            rom[14077] = 8'hf3 ;
            rom[14078] = 8'hec ;
            rom[14079] = 8'hde ;
            rom[14080] = 8'h0b ;
            rom[14081] = 8'hfa ;
            rom[14082] = 8'hef ;
            rom[14083] = 8'hee ;
            rom[14084] = 8'h0b ;
            rom[14085] = 8'he1 ;
            rom[14086] = 8'h03 ;
            rom[14087] = 8'hf3 ;
            rom[14088] = 8'hd6 ;
            rom[14089] = 8'h39 ;
            rom[14090] = 8'hf6 ;
            rom[14091] = 8'hf6 ;
            rom[14092] = 8'h03 ;
            rom[14093] = 8'h0d ;
            rom[14094] = 8'hea ;
            rom[14095] = 8'hed ;
            rom[14096] = 8'hf4 ;
            rom[14097] = 8'he8 ;
            rom[14098] = 8'h1f ;
            rom[14099] = 8'hd6 ;
            rom[14100] = 8'he5 ;
            rom[14101] = 8'he0 ;
            rom[14102] = 8'heb ;
            rom[14103] = 8'hee ;
            rom[14104] = 8'h9c ;
            rom[14105] = 8'h20 ;
            rom[14106] = 8'hfd ;
            rom[14107] = 8'hf0 ;
            rom[14108] = 8'h17 ;
            rom[14109] = 8'h06 ;
            rom[14110] = 8'h17 ;
            rom[14111] = 8'h00 ;
            rom[14112] = 8'hf7 ;
            rom[14113] = 8'he1 ;
            rom[14114] = 8'h1a ;
            rom[14115] = 8'hed ;
            rom[14116] = 8'he6 ;
            rom[14117] = 8'hf0 ;
            rom[14118] = 8'h03 ;
            rom[14119] = 8'hfd ;
            rom[14120] = 8'h1d ;
            rom[14121] = 8'h1b ;
            rom[14122] = 8'hed ;
            rom[14123] = 8'hbb ;
            rom[14124] = 8'hf0 ;
            rom[14125] = 8'hf6 ;
            rom[14126] = 8'h06 ;
            rom[14127] = 8'hd2 ;
            rom[14128] = 8'h0d ;
            rom[14129] = 8'he1 ;
            rom[14130] = 8'hdd ;
            rom[14131] = 8'hee ;
            rom[14132] = 8'heb ;
            rom[14133] = 8'hf5 ;
            rom[14134] = 8'hef ;
            rom[14135] = 8'hf5 ;
            rom[14136] = 8'hcc ;
            rom[14137] = 8'hfc ;
            rom[14138] = 8'h1c ;
            rom[14139] = 8'h2b ;
            rom[14140] = 8'h17 ;
            rom[14141] = 8'hfe ;
            rom[14142] = 8'hec ;
            rom[14143] = 8'h2d ;
            rom[14144] = 8'he1 ;
            rom[14145] = 8'hfe ;
            rom[14146] = 8'h02 ;
            rom[14147] = 8'hcf ;
            rom[14148] = 8'h04 ;
            rom[14149] = 8'h09 ;
            rom[14150] = 8'hd9 ;
            rom[14151] = 8'h15 ;
            rom[14152] = 8'hfe ;
            rom[14153] = 8'h16 ;
            rom[14154] = 8'h0e ;
            rom[14155] = 8'h15 ;
            rom[14156] = 8'hd5 ;
            rom[14157] = 8'he9 ;
            rom[14158] = 8'hf1 ;
            rom[14159] = 8'hfe ;
            rom[14160] = 8'he9 ;
            rom[14161] = 8'he4 ;
            rom[14162] = 8'hda ;
            rom[14163] = 8'hf9 ;
            rom[14164] = 8'h17 ;
            rom[14165] = 8'hf0 ;
            rom[14166] = 8'hf2 ;
            rom[14167] = 8'h2d ;
            rom[14168] = 8'he5 ;
            rom[14169] = 8'hc9 ;
            rom[14170] = 8'hdc ;
            rom[14171] = 8'hd5 ;
            rom[14172] = 8'he5 ;
            rom[14173] = 8'he0 ;
            rom[14174] = 8'hf9 ;
            rom[14175] = 8'h1c ;
            rom[14176] = 8'hf1 ;
            rom[14177] = 8'hc5 ;
            rom[14178] = 8'hd3 ;
            rom[14179] = 8'hf0 ;
            rom[14180] = 8'hfb ;
            rom[14181] = 8'h07 ;
            rom[14182] = 8'h05 ;
            rom[14183] = 8'heb ;
            rom[14184] = 8'he1 ;
            rom[14185] = 8'hfc ;
            rom[14186] = 8'h0b ;
            rom[14187] = 8'he4 ;
            rom[14188] = 8'he8 ;
            rom[14189] = 8'hca ;
            rom[14190] = 8'h12 ;
            rom[14191] = 8'hda ;
            rom[14192] = 8'hd0 ;
            rom[14193] = 8'he6 ;
            rom[14194] = 8'h18 ;
            rom[14195] = 8'he3 ;
            rom[14196] = 8'h1e ;
            rom[14197] = 8'h0f ;
            rom[14198] = 8'h0d ;
            rom[14199] = 8'hcf ;
            rom[14200] = 8'hdd ;
            rom[14201] = 8'h0c ;
            rom[14202] = 8'h0f ;
            rom[14203] = 8'hfa ;
            rom[14204] = 8'h29 ;
            rom[14205] = 8'hdb ;
            rom[14206] = 8'hfd ;
            rom[14207] = 8'hcd ;
            rom[14208] = 8'hcd ;
            rom[14209] = 8'h03 ;
            rom[14210] = 8'hea ;
            rom[14211] = 8'heb ;
            rom[14212] = 8'hf4 ;
            rom[14213] = 8'he1 ;
            rom[14214] = 8'hcf ;
            rom[14215] = 8'h1c ;
            rom[14216] = 8'hf3 ;
            rom[14217] = 8'hfa ;
            rom[14218] = 8'hd0 ;
            rom[14219] = 8'h01 ;
            rom[14220] = 8'hec ;
            rom[14221] = 8'h01 ;
            rom[14222] = 8'h19 ;
            rom[14223] = 8'hf7 ;
            rom[14224] = 8'h0c ;
            rom[14225] = 8'hf9 ;
            rom[14226] = 8'hf1 ;
            rom[14227] = 8'hf3 ;
            rom[14228] = 8'hec ;
            rom[14229] = 8'hff ;
            rom[14230] = 8'h06 ;
            rom[14231] = 8'h1c ;
            rom[14232] = 8'h1b ;
            rom[14233] = 8'he4 ;
            rom[14234] = 8'hfe ;
            rom[14235] = 8'he8 ;
            rom[14236] = 8'hcb ;
            rom[14237] = 8'h09 ;
            rom[14238] = 8'h13 ;
            rom[14239] = 8'h10 ;
            rom[14240] = 8'h27 ;
            rom[14241] = 8'h0b ;
            rom[14242] = 8'h16 ;
            rom[14243] = 8'he8 ;
            rom[14244] = 8'hf1 ;
            rom[14245] = 8'hf5 ;
            rom[14246] = 8'h02 ;
            rom[14247] = 8'hda ;
            rom[14248] = 8'hde ;
            rom[14249] = 8'hc7 ;
            rom[14250] = 8'hd9 ;
            rom[14251] = 8'h0f ;
            rom[14252] = 8'h17 ;
            rom[14253] = 8'hee ;
            rom[14254] = 8'hbd ;
            rom[14255] = 8'hfe ;
            rom[14256] = 8'h0a ;
            rom[14257] = 8'hdc ;
            rom[14258] = 8'h07 ;
            rom[14259] = 8'hec ;
            rom[14260] = 8'hf8 ;
            rom[14261] = 8'hf9 ;
            rom[14262] = 8'h0f ;
            rom[14263] = 8'h08 ;
            rom[14264] = 8'h00 ;
            rom[14265] = 8'hfa ;
            rom[14266] = 8'h0e ;
            rom[14267] = 8'hf5 ;
            rom[14268] = 8'h03 ;
            rom[14269] = 8'hdc ;
            rom[14270] = 8'h0d ;
            rom[14271] = 8'h0f ;
            rom[14272] = 8'h1f ;
            rom[14273] = 8'hf3 ;
            rom[14274] = 8'h12 ;
            rom[14275] = 8'hf8 ;
            rom[14276] = 8'h0f ;
            rom[14277] = 8'h0a ;
            rom[14278] = 8'hea ;
            rom[14279] = 8'hd7 ;
            rom[14280] = 8'hee ;
            rom[14281] = 8'hf7 ;
            rom[14282] = 8'hfb ;
            rom[14283] = 8'hf8 ;
            rom[14284] = 8'h15 ;
            rom[14285] = 8'he6 ;
            rom[14286] = 8'hf1 ;
            rom[14287] = 8'h08 ;
            rom[14288] = 8'h05 ;
            rom[14289] = 8'h14 ;
            rom[14290] = 8'h39 ;
            rom[14291] = 8'he1 ;
            rom[14292] = 8'hfc ;
            rom[14293] = 8'hff ;
            rom[14294] = 8'hba ;
            rom[14295] = 8'hec ;
            rom[14296] = 8'hdf ;
            rom[14297] = 8'h0d ;
            rom[14298] = 8'hf0 ;
            rom[14299] = 8'h12 ;
            rom[14300] = 8'hfe ;
            rom[14301] = 8'h21 ;
            rom[14302] = 8'h04 ;
            rom[14303] = 8'hf4 ;
            rom[14304] = 8'h14 ;
            rom[14305] = 8'h06 ;
            rom[14306] = 8'h0a ;
            rom[14307] = 8'hf6 ;
            rom[14308] = 8'hf0 ;
            rom[14309] = 8'h10 ;
            rom[14310] = 8'h0a ;
            rom[14311] = 8'hef ;
            rom[14312] = 8'h18 ;
            rom[14313] = 8'h2b ;
            rom[14314] = 8'hf7 ;
            rom[14315] = 8'h2a ;
            rom[14316] = 8'hfe ;
            rom[14317] = 8'h05 ;
            rom[14318] = 8'heb ;
            rom[14319] = 8'hf1 ;
            rom[14320] = 8'h11 ;
            rom[14321] = 8'h11 ;
            rom[14322] = 8'heb ;
            rom[14323] = 8'hfa ;
            rom[14324] = 8'h09 ;
            rom[14325] = 8'hfe ;
            rom[14326] = 8'hf6 ;
            rom[14327] = 8'h0e ;
            rom[14328] = 8'hd8 ;
            rom[14329] = 8'h10 ;
            rom[14330] = 8'he8 ;
            rom[14331] = 8'he9 ;
            rom[14332] = 8'hde ;
            rom[14333] = 8'h2f ;
            rom[14334] = 8'h16 ;
            rom[14335] = 8'h2e ;
            rom[14336] = 8'hdc ;
            rom[14337] = 8'he3 ;
            rom[14338] = 8'hdb ;
            rom[14339] = 8'hfa ;
            rom[14340] = 8'h0e ;
            rom[14341] = 8'h09 ;
            rom[14342] = 8'hf5 ;
            rom[14343] = 8'h01 ;
            rom[14344] = 8'h05 ;
            rom[14345] = 8'he2 ;
            rom[14346] = 8'he3 ;
            rom[14347] = 8'hea ;
            rom[14348] = 8'hf2 ;
            rom[14349] = 8'hea ;
            rom[14350] = 8'h1c ;
            rom[14351] = 8'h07 ;
            rom[14352] = 8'h0c ;
            rom[14353] = 8'he8 ;
            rom[14354] = 8'hd6 ;
            rom[14355] = 8'h07 ;
            rom[14356] = 8'hf9 ;
            rom[14357] = 8'heb ;
            rom[14358] = 8'h17 ;
            rom[14359] = 8'h0b ;
            rom[14360] = 8'h08 ;
            rom[14361] = 8'hfe ;
            rom[14362] = 8'h1e ;
            rom[14363] = 8'hfb ;
            rom[14364] = 8'hf9 ;
            rom[14365] = 8'h09 ;
            rom[14366] = 8'hd4 ;
            rom[14367] = 8'h04 ;
            rom[14368] = 8'h25 ;
            rom[14369] = 8'hf5 ;
            rom[14370] = 8'hd9 ;
            rom[14371] = 8'hfd ;
            rom[14372] = 8'hf8 ;
            rom[14373] = 8'hf5 ;
            rom[14374] = 8'hfb ;
            rom[14375] = 8'h18 ;
            rom[14376] = 8'h12 ;
            rom[14377] = 8'hfc ;
            rom[14378] = 8'h01 ;
            rom[14379] = 8'hd9 ;
            rom[14380] = 8'hda ;
            rom[14381] = 8'h0a ;
            rom[14382] = 8'hd7 ;
            rom[14383] = 8'h03 ;
            rom[14384] = 8'h0b ;
            rom[14385] = 8'he9 ;
            rom[14386] = 8'h07 ;
            rom[14387] = 8'heb ;
            rom[14388] = 8'h11 ;
            rom[14389] = 8'hf7 ;
            rom[14390] = 8'hfe ;
            rom[14391] = 8'h1e ;
            rom[14392] = 8'heb ;
            rom[14393] = 8'h00 ;
            rom[14394] = 8'h09 ;
            rom[14395] = 8'hec ;
            rom[14396] = 8'hf9 ;
            rom[14397] = 8'hd9 ;
            rom[14398] = 8'he6 ;
            rom[14399] = 8'hf7 ;
            rom[14400] = 8'hff ;
            rom[14401] = 8'he2 ;
            rom[14402] = 8'h10 ;
            rom[14403] = 8'h0a ;
            rom[14404] = 8'h01 ;
            rom[14405] = 8'h15 ;
            rom[14406] = 8'hff ;
            rom[14407] = 8'hf0 ;
            rom[14408] = 8'h1c ;
            rom[14409] = 8'hcd ;
            rom[14410] = 8'hff ;
            rom[14411] = 8'hfa ;
            rom[14412] = 8'h00 ;
            rom[14413] = 8'hdd ;
            rom[14414] = 8'hfa ;
            rom[14415] = 8'h13 ;
            rom[14416] = 8'he4 ;
            rom[14417] = 8'he4 ;
            rom[14418] = 8'h12 ;
            rom[14419] = 8'hed ;
            rom[14420] = 8'hdf ;
            rom[14421] = 8'h17 ;
            rom[14422] = 8'hdf ;
            rom[14423] = 8'hf9 ;
            rom[14424] = 8'he2 ;
            rom[14425] = 8'h0b ;
            rom[14426] = 8'hf1 ;
            rom[14427] = 8'h00 ;
            rom[14428] = 8'hff ;
            rom[14429] = 8'heb ;
            rom[14430] = 8'h04 ;
            rom[14431] = 8'hf5 ;
            rom[14432] = 8'h04 ;
            rom[14433] = 8'hfe ;
            rom[14434] = 8'h01 ;
            rom[14435] = 8'hcf ;
            rom[14436] = 8'he4 ;
            rom[14437] = 8'he5 ;
            rom[14438] = 8'h05 ;
            rom[14439] = 8'h04 ;
            rom[14440] = 8'h13 ;
            rom[14441] = 8'hf1 ;
            rom[14442] = 8'hd4 ;
            rom[14443] = 8'h0f ;
            rom[14444] = 8'h33 ;
            rom[14445] = 8'h19 ;
            rom[14446] = 8'hdb ;
            rom[14447] = 8'h13 ;
            rom[14448] = 8'hf9 ;
            rom[14449] = 8'hfa ;
            rom[14450] = 8'h13 ;
            rom[14451] = 8'h07 ;
            rom[14452] = 8'he3 ;
            rom[14453] = 8'he4 ;
            rom[14454] = 8'h1c ;
            rom[14455] = 8'h12 ;
            rom[14456] = 8'hff ;
            rom[14457] = 8'hfc ;
            rom[14458] = 8'hf5 ;
            rom[14459] = 8'hf0 ;
            rom[14460] = 8'hed ;
            rom[14461] = 8'h0e ;
            rom[14462] = 8'h12 ;
            rom[14463] = 8'hf7 ;
            rom[14464] = 8'he6 ;
            rom[14465] = 8'ha5 ;
            rom[14466] = 8'h09 ;
            rom[14467] = 8'h24 ;
            rom[14468] = 8'hda ;
            rom[14469] = 8'h02 ;
            rom[14470] = 8'hcf ;
            rom[14471] = 8'h11 ;
            rom[14472] = 8'h00 ;
            rom[14473] = 8'hd9 ;
            rom[14474] = 8'h16 ;
            rom[14475] = 8'hfb ;
            rom[14476] = 8'h22 ;
            rom[14477] = 8'hf3 ;
            rom[14478] = 8'h27 ;
            rom[14479] = 8'he9 ;
            rom[14480] = 8'h0e ;
            rom[14481] = 8'h18 ;
            rom[14482] = 8'hdf ;
            rom[14483] = 8'h26 ;
            rom[14484] = 8'h1d ;
            rom[14485] = 8'h17 ;
            rom[14486] = 8'hfe ;
            rom[14487] = 8'hf8 ;
            rom[14488] = 8'h33 ;
            rom[14489] = 8'h05 ;
            rom[14490] = 8'hfd ;
            rom[14491] = 8'he6 ;
            rom[14492] = 8'hd2 ;
            rom[14493] = 8'h01 ;
            rom[14494] = 8'h00 ;
            rom[14495] = 8'h13 ;
            rom[14496] = 8'hfe ;
            rom[14497] = 8'h01 ;
            rom[14498] = 8'hfd ;
            rom[14499] = 8'he6 ;
            rom[14500] = 8'h03 ;
            rom[14501] = 8'h00 ;
            rom[14502] = 8'h09 ;
            rom[14503] = 8'hf0 ;
            rom[14504] = 8'hf9 ;
            rom[14505] = 8'hf5 ;
            rom[14506] = 8'he2 ;
            rom[14507] = 8'hf5 ;
            rom[14508] = 8'hf1 ;
            rom[14509] = 8'h0a ;
            rom[14510] = 8'hca ;
            rom[14511] = 8'hfd ;
            rom[14512] = 8'he5 ;
            rom[14513] = 8'hf7 ;
            rom[14514] = 8'hfc ;
            rom[14515] = 8'h03 ;
            rom[14516] = 8'h03 ;
            rom[14517] = 8'hd8 ;
            rom[14518] = 8'heb ;
            rom[14519] = 8'h02 ;
            rom[14520] = 8'hef ;
            rom[14521] = 8'he8 ;
            rom[14522] = 8'h19 ;
            rom[14523] = 8'he1 ;
            rom[14524] = 8'hfb ;
            rom[14525] = 8'hd1 ;
            rom[14526] = 8'he6 ;
            rom[14527] = 8'hf3 ;
            rom[14528] = 8'hd9 ;
            rom[14529] = 8'hf9 ;
            rom[14530] = 8'hfa ;
            rom[14531] = 8'hed ;
            rom[14532] = 8'h21 ;
            rom[14533] = 8'hed ;
            rom[14534] = 8'h06 ;
            rom[14535] = 8'hfa ;
            rom[14536] = 8'h1b ;
            rom[14537] = 8'h0d ;
            rom[14538] = 8'hf9 ;
            rom[14539] = 8'h0c ;
            rom[14540] = 8'hd9 ;
            rom[14541] = 8'h01 ;
            rom[14542] = 8'hfc ;
            rom[14543] = 8'hed ;
            rom[14544] = 8'he7 ;
            rom[14545] = 8'hf0 ;
            rom[14546] = 8'h11 ;
            rom[14547] = 8'hcb ;
            rom[14548] = 8'h1c ;
            rom[14549] = 8'h1d ;
            rom[14550] = 8'h05 ;
            rom[14551] = 8'he5 ;
            rom[14552] = 8'hd7 ;
            rom[14553] = 8'he9 ;
            rom[14554] = 8'h0e ;
            rom[14555] = 8'h24 ;
            rom[14556] = 8'h1d ;
            rom[14557] = 8'hdb ;
            rom[14558] = 8'hfc ;
            rom[14559] = 8'hea ;
            rom[14560] = 8'h06 ;
            rom[14561] = 8'hfb ;
            rom[14562] = 8'hf7 ;
            rom[14563] = 8'h08 ;
            rom[14564] = 8'hea ;
            rom[14565] = 8'h31 ;
            rom[14566] = 8'hfc ;
            rom[14567] = 8'hfb ;
            rom[14568] = 8'hf9 ;
            rom[14569] = 8'hf2 ;
            rom[14570] = 8'h0b ;
            rom[14571] = 8'hff ;
            rom[14572] = 8'h2d ;
            rom[14573] = 8'h13 ;
            rom[14574] = 8'h23 ;
            rom[14575] = 8'hea ;
            rom[14576] = 8'hda ;
            rom[14577] = 8'hfb ;
            rom[14578] = 8'h18 ;
            rom[14579] = 8'hba ;
            rom[14580] = 8'hf7 ;
            rom[14581] = 8'hee ;
            rom[14582] = 8'he9 ;
            rom[14583] = 8'h11 ;
            rom[14584] = 8'hec ;
            rom[14585] = 8'hf5 ;
            rom[14586] = 8'h1e ;
            rom[14587] = 8'hf3 ;
            rom[14588] = 8'hc1 ;
            rom[14589] = 8'hf3 ;
            rom[14590] = 8'hf9 ;
            rom[14591] = 8'h25 ;
            rom[14592] = 8'h06 ;
            rom[14593] = 8'h0e ;
            rom[14594] = 8'hfc ;
            rom[14595] = 8'hfc ;
            rom[14596] = 8'hf9 ;
            rom[14597] = 8'hf6 ;
            rom[14598] = 8'h16 ;
            rom[14599] = 8'he0 ;
            rom[14600] = 8'hd8 ;
            rom[14601] = 8'hcc ;
            rom[14602] = 8'hd9 ;
            rom[14603] = 8'hfb ;
            rom[14604] = 8'hdd ;
            rom[14605] = 8'he4 ;
            rom[14606] = 8'h00 ;
            rom[14607] = 8'h24 ;
            rom[14608] = 8'hfc ;
            rom[14609] = 8'h07 ;
            rom[14610] = 8'h19 ;
            rom[14611] = 8'hfb ;
            rom[14612] = 8'hee ;
            rom[14613] = 8'hf2 ;
            rom[14614] = 8'hf0 ;
            rom[14615] = 8'h19 ;
            rom[14616] = 8'hd2 ;
            rom[14617] = 8'hf1 ;
            rom[14618] = 8'heb ;
            rom[14619] = 8'hf3 ;
            rom[14620] = 8'hfd ;
            rom[14621] = 8'h2a ;
            rom[14622] = 8'h18 ;
            rom[14623] = 8'hf0 ;
            rom[14624] = 8'hc9 ;
            rom[14625] = 8'hf4 ;
            rom[14626] = 8'hfd ;
            rom[14627] = 8'hf4 ;
            rom[14628] = 8'hd0 ;
            rom[14629] = 8'hfe ;
            rom[14630] = 8'h04 ;
            rom[14631] = 8'h06 ;
            rom[14632] = 8'h11 ;
            rom[14633] = 8'h12 ;
            rom[14634] = 8'h08 ;
            rom[14635] = 8'h22 ;
            rom[14636] = 8'h22 ;
            rom[14637] = 8'h00 ;
            rom[14638] = 8'hfb ;
            rom[14639] = 8'hf6 ;
            rom[14640] = 8'hc8 ;
            rom[14641] = 8'hc7 ;
            rom[14642] = 8'h11 ;
            rom[14643] = 8'hfe ;
            rom[14644] = 8'he4 ;
            rom[14645] = 8'hfa ;
            rom[14646] = 8'hf3 ;
            rom[14647] = 8'h01 ;
            rom[14648] = 8'h0b ;
            rom[14649] = 8'hf5 ;
            rom[14650] = 8'h12 ;
            rom[14651] = 8'hd4 ;
            rom[14652] = 8'h23 ;
            rom[14653] = 8'hdc ;
            rom[14654] = 8'h14 ;
            rom[14655] = 8'h06 ;
            rom[14656] = 8'he5 ;
            rom[14657] = 8'h16 ;
            rom[14658] = 8'hce ;
            rom[14659] = 8'h17 ;
            rom[14660] = 8'hc1 ;
            rom[14661] = 8'h0f ;
            rom[14662] = 8'hcf ;
            rom[14663] = 8'h02 ;
            rom[14664] = 8'hd2 ;
            rom[14665] = 8'h16 ;
            rom[14666] = 8'hfd ;
            rom[14667] = 8'hdc ;
            rom[14668] = 8'h10 ;
            rom[14669] = 8'h04 ;
            rom[14670] = 8'hfa ;
            rom[14671] = 8'h00 ;
            rom[14672] = 8'hfa ;
            rom[14673] = 8'h0a ;
            rom[14674] = 8'h0f ;
            rom[14675] = 8'h06 ;
            rom[14676] = 8'h04 ;
            rom[14677] = 8'h0a ;
            rom[14678] = 8'hf7 ;
            rom[14679] = 8'h39 ;
            rom[14680] = 8'he6 ;
            rom[14681] = 8'h17 ;
            rom[14682] = 8'h04 ;
            rom[14683] = 8'hfc ;
            rom[14684] = 8'hfd ;
            rom[14685] = 8'hcc ;
            rom[14686] = 8'h0f ;
            rom[14687] = 8'h0c ;
            rom[14688] = 8'h1e ;
            rom[14689] = 8'h15 ;
            rom[14690] = 8'heb ;
            rom[14691] = 8'hee ;
            rom[14692] = 8'he7 ;
            rom[14693] = 8'hf2 ;
            rom[14694] = 8'hf1 ;
            rom[14695] = 8'hf8 ;
            rom[14696] = 8'h08 ;
            rom[14697] = 8'h0f ;
            rom[14698] = 8'hf1 ;
            rom[14699] = 8'h0a ;
            rom[14700] = 8'hcf ;
            rom[14701] = 8'hd8 ;
            rom[14702] = 8'h14 ;
            rom[14703] = 8'h01 ;
            rom[14704] = 8'h05 ;
            rom[14705] = 8'he9 ;
            rom[14706] = 8'h02 ;
            rom[14707] = 8'h4b ;
            rom[14708] = 8'h25 ;
            rom[14709] = 8'h17 ;
            rom[14710] = 8'hff ;
            rom[14711] = 8'h0d ;
            rom[14712] = 8'h00 ;
            rom[14713] = 8'h08 ;
            rom[14714] = 8'hec ;
            rom[14715] = 8'heb ;
            rom[14716] = 8'h18 ;
            rom[14717] = 8'h10 ;
            rom[14718] = 8'h1b ;
            rom[14719] = 8'h05 ;
            rom[14720] = 8'hfa ;
            rom[14721] = 8'he0 ;
            rom[14722] = 8'hfc ;
            rom[14723] = 8'hdc ;
            rom[14724] = 8'h05 ;
            rom[14725] = 8'h13 ;
            rom[14726] = 8'hfe ;
            rom[14727] = 8'h0e ;
            rom[14728] = 8'h1d ;
            rom[14729] = 8'he2 ;
            rom[14730] = 8'h29 ;
            rom[14731] = 8'hf5 ;
            rom[14732] = 8'h09 ;
            rom[14733] = 8'h0d ;
            rom[14734] = 8'h0c ;
            rom[14735] = 8'hcf ;
            rom[14736] = 8'hd5 ;
            rom[14737] = 8'h0f ;
            rom[14738] = 8'hfc ;
            rom[14739] = 8'h10 ;
            rom[14740] = 8'hcb ;
            rom[14741] = 8'hf1 ;
            rom[14742] = 8'h07 ;
            rom[14743] = 8'h20 ;
            rom[14744] = 8'h19 ;
            rom[14745] = 8'hf9 ;
            rom[14746] = 8'hc5 ;
            rom[14747] = 8'hfa ;
            rom[14748] = 8'h22 ;
            rom[14749] = 8'h0d ;
            rom[14750] = 8'h00 ;
            rom[14751] = 8'hf5 ;
            rom[14752] = 8'hd6 ;
            rom[14753] = 8'he9 ;
            rom[14754] = 8'h19 ;
            rom[14755] = 8'hf2 ;
            rom[14756] = 8'h16 ;
            rom[14757] = 8'hea ;
            rom[14758] = 8'h10 ;
            rom[14759] = 8'hf5 ;
            rom[14760] = 8'h05 ;
            rom[14761] = 8'hed ;
            rom[14762] = 8'hf9 ;
            rom[14763] = 8'h1a ;
            rom[14764] = 8'h10 ;
            rom[14765] = 8'h01 ;
            rom[14766] = 8'h19 ;
            rom[14767] = 8'hd1 ;
            rom[14768] = 8'h20 ;
            rom[14769] = 8'hfa ;
            rom[14770] = 8'hd2 ;
            rom[14771] = 8'h15 ;
            rom[14772] = 8'h0b ;
            rom[14773] = 8'hf0 ;
            rom[14774] = 8'hfe ;
            rom[14775] = 8'h1a ;
            rom[14776] = 8'h08 ;
            rom[14777] = 8'h05 ;
            rom[14778] = 8'h00 ;
            rom[14779] = 8'h18 ;
            rom[14780] = 8'h16 ;
            rom[14781] = 8'hca ;
            rom[14782] = 8'h0c ;
            rom[14783] = 8'hfb ;
            rom[14784] = 8'h0d ;
            rom[14785] = 8'h14 ;
            rom[14786] = 8'h0f ;
            rom[14787] = 8'he5 ;
            rom[14788] = 8'h04 ;
            rom[14789] = 8'h13 ;
            rom[14790] = 8'h0c ;
            rom[14791] = 8'he4 ;
            rom[14792] = 8'hfe ;
            rom[14793] = 8'hf6 ;
            rom[14794] = 8'hf9 ;
            rom[14795] = 8'hfb ;
            rom[14796] = 8'he0 ;
            rom[14797] = 8'h08 ;
            rom[14798] = 8'h10 ;
            rom[14799] = 8'he9 ;
            rom[14800] = 8'h05 ;
            rom[14801] = 8'hfd ;
            rom[14802] = 8'he7 ;
            rom[14803] = 8'h03 ;
            rom[14804] = 8'hde ;
            rom[14805] = 8'h15 ;
            rom[14806] = 8'he0 ;
            rom[14807] = 8'heb ;
            rom[14808] = 8'hef ;
            rom[14809] = 8'h08 ;
            rom[14810] = 8'hec ;
            rom[14811] = 8'h0a ;
            rom[14812] = 8'h07 ;
            rom[14813] = 8'h14 ;
            rom[14814] = 8'hd7 ;
            rom[14815] = 8'hfb ;
            rom[14816] = 8'h04 ;
            rom[14817] = 8'hea ;
            rom[14818] = 8'hf3 ;
            rom[14819] = 8'h06 ;
            rom[14820] = 8'h0a ;
            rom[14821] = 8'hf7 ;
            rom[14822] = 8'hff ;
            rom[14823] = 8'h15 ;
            rom[14824] = 8'hf6 ;
            rom[14825] = 8'hfa ;
            rom[14826] = 8'h28 ;
            rom[14827] = 8'hfd ;
            rom[14828] = 8'h23 ;
            rom[14829] = 8'hb7 ;
            rom[14830] = 8'h17 ;
            rom[14831] = 8'he9 ;
            rom[14832] = 8'he5 ;
            rom[14833] = 8'hee ;
            rom[14834] = 8'h2e ;
            rom[14835] = 8'h03 ;
            rom[14836] = 8'h11 ;
            rom[14837] = 8'hdc ;
            rom[14838] = 8'h0f ;
            rom[14839] = 8'hf1 ;
            rom[14840] = 8'hed ;
            rom[14841] = 8'h0b ;
            rom[14842] = 8'h18 ;
            rom[14843] = 8'h18 ;
            rom[14844] = 8'hea ;
            rom[14845] = 8'hfd ;
            rom[14846] = 8'h15 ;
            rom[14847] = 8'h09 ;
            rom[14848] = 8'he7 ;
            rom[14849] = 8'hf9 ;
            rom[14850] = 8'hee ;
            rom[14851] = 8'h07 ;
            rom[14852] = 8'h07 ;
            rom[14853] = 8'hfe ;
            rom[14854] = 8'hfe ;
            rom[14855] = 8'hf6 ;
            rom[14856] = 8'hd7 ;
            rom[14857] = 8'hee ;
            rom[14858] = 8'h17 ;
            rom[14859] = 8'h16 ;
            rom[14860] = 8'hf7 ;
            rom[14861] = 8'hc4 ;
            rom[14862] = 8'hef ;
            rom[14863] = 8'hf8 ;
            rom[14864] = 8'hf9 ;
            rom[14865] = 8'hca ;
            rom[14866] = 8'h0c ;
            rom[14867] = 8'he4 ;
            rom[14868] = 8'h05 ;
            rom[14869] = 8'h02 ;
            rom[14870] = 8'h09 ;
            rom[14871] = 8'hd1 ;
            rom[14872] = 8'h05 ;
            rom[14873] = 8'he8 ;
            rom[14874] = 8'hf1 ;
            rom[14875] = 8'hf4 ;
            rom[14876] = 8'h14 ;
            rom[14877] = 8'h06 ;
            rom[14878] = 8'hf9 ;
            rom[14879] = 8'hf8 ;
            rom[14880] = 8'h25 ;
            rom[14881] = 8'hf8 ;
            rom[14882] = 8'hf9 ;
            rom[14883] = 8'h19 ;
            rom[14884] = 8'h12 ;
            rom[14885] = 8'h01 ;
            rom[14886] = 8'h02 ;
            rom[14887] = 8'h22 ;
            rom[14888] = 8'hf3 ;
            rom[14889] = 8'hee ;
            rom[14890] = 8'hfd ;
            rom[14891] = 8'he2 ;
            rom[14892] = 8'hf3 ;
            rom[14893] = 8'h0b ;
            rom[14894] = 8'hf3 ;
            rom[14895] = 8'h16 ;
            rom[14896] = 8'h19 ;
            rom[14897] = 8'hf6 ;
            rom[14898] = 8'hfe ;
            rom[14899] = 8'h05 ;
            rom[14900] = 8'hdd ;
            rom[14901] = 8'h0a ;
            rom[14902] = 8'hd2 ;
            rom[14903] = 8'hde ;
            rom[14904] = 8'hfc ;
            rom[14905] = 8'h1d ;
            rom[14906] = 8'hea ;
            rom[14907] = 8'h0c ;
            rom[14908] = 8'h17 ;
            rom[14909] = 8'h02 ;
            rom[14910] = 8'h06 ;
            rom[14911] = 8'hd5 ;
            rom[14912] = 8'hf8 ;
            rom[14913] = 8'h14 ;
            rom[14914] = 8'hfb ;
            rom[14915] = 8'hfc ;
            rom[14916] = 8'hd2 ;
            rom[14917] = 8'h26 ;
            rom[14918] = 8'h08 ;
            rom[14919] = 8'h11 ;
            rom[14920] = 8'hec ;
            rom[14921] = 8'he0 ;
            rom[14922] = 8'h11 ;
            rom[14923] = 8'hfc ;
            rom[14924] = 8'he5 ;
            rom[14925] = 8'hf4 ;
            rom[14926] = 8'hdd ;
            rom[14927] = 8'hf2 ;
            rom[14928] = 8'h2d ;
            rom[14929] = 8'he5 ;
            rom[14930] = 8'h04 ;
            rom[14931] = 8'hdc ;
            rom[14932] = 8'hf0 ;
            rom[14933] = 8'he3 ;
            rom[14934] = 8'h24 ;
            rom[14935] = 8'hf6 ;
            rom[14936] = 8'h06 ;
            rom[14937] = 8'hf9 ;
            rom[14938] = 8'h10 ;
            rom[14939] = 8'h0c ;
            rom[14940] = 8'hfa ;
            rom[14941] = 8'he2 ;
            rom[14942] = 8'hdd ;
            rom[14943] = 8'hf8 ;
            rom[14944] = 8'hea ;
            rom[14945] = 8'h19 ;
            rom[14946] = 8'he9 ;
            rom[14947] = 8'hbb ;
            rom[14948] = 8'hf4 ;
            rom[14949] = 8'h29 ;
            rom[14950] = 8'h2e ;
            rom[14951] = 8'h28 ;
            rom[14952] = 8'hf0 ;
            rom[14953] = 8'h06 ;
            rom[14954] = 8'h22 ;
            rom[14955] = 8'hfe ;
            rom[14956] = 8'hf5 ;
            rom[14957] = 8'hec ;
            rom[14958] = 8'hf0 ;
            rom[14959] = 8'h0e ;
            rom[14960] = 8'hf7 ;
            rom[14961] = 8'hf5 ;
            rom[14962] = 8'h1a ;
            rom[14963] = 8'h05 ;
            rom[14964] = 8'hee ;
            rom[14965] = 8'h17 ;
            rom[14966] = 8'hf3 ;
            rom[14967] = 8'hfa ;
            rom[14968] = 8'hf0 ;
            rom[14969] = 8'hfd ;
            rom[14970] = 8'h10 ;
            rom[14971] = 8'hec ;
            rom[14972] = 8'hd5 ;
            rom[14973] = 8'h05 ;
            rom[14974] = 8'h07 ;
            rom[14975] = 8'hf6 ;
            rom[14976] = 8'he6 ;
            rom[14977] = 8'h06 ;
            rom[14978] = 8'hfd ;
            rom[14979] = 8'h28 ;
            rom[14980] = 8'h0a ;
            rom[14981] = 8'h0a ;
            rom[14982] = 8'he8 ;
            rom[14983] = 8'h1b ;
            rom[14984] = 8'h26 ;
            rom[14985] = 8'he2 ;
            rom[14986] = 8'hef ;
            rom[14987] = 8'hf7 ;
            rom[14988] = 8'hd9 ;
            rom[14989] = 8'h17 ;
            rom[14990] = 8'h13 ;
            rom[14991] = 8'hf6 ;
            rom[14992] = 8'h09 ;
            rom[14993] = 8'h0b ;
            rom[14994] = 8'he9 ;
            rom[14995] = 8'hd5 ;
            rom[14996] = 8'h05 ;
            rom[14997] = 8'h0f ;
            rom[14998] = 8'h0e ;
            rom[14999] = 8'h0d ;
            rom[15000] = 8'h14 ;
            rom[15001] = 8'he7 ;
            rom[15002] = 8'h1b ;
            rom[15003] = 8'h15 ;
            rom[15004] = 8'hf5 ;
            rom[15005] = 8'hfe ;
            rom[15006] = 8'h08 ;
            rom[15007] = 8'h0e ;
            rom[15008] = 8'h2a ;
            rom[15009] = 8'hf2 ;
            rom[15010] = 8'h14 ;
            rom[15011] = 8'hd4 ;
            rom[15012] = 8'hdb ;
            rom[15013] = 8'hf9 ;
            rom[15014] = 8'h23 ;
            rom[15015] = 8'h0b ;
            rom[15016] = 8'hf9 ;
            rom[15017] = 8'hf4 ;
            rom[15018] = 8'hff ;
            rom[15019] = 8'h1b ;
            rom[15020] = 8'h31 ;
            rom[15021] = 8'hf7 ;
            rom[15022] = 8'hfd ;
            rom[15023] = 8'h0f ;
            rom[15024] = 8'he2 ;
            rom[15025] = 8'h00 ;
            rom[15026] = 8'hf2 ;
            rom[15027] = 8'hdb ;
            rom[15028] = 8'h11 ;
            rom[15029] = 8'he8 ;
            rom[15030] = 8'h00 ;
            rom[15031] = 8'hef ;
            rom[15032] = 8'h12 ;
            rom[15033] = 8'hf2 ;
            rom[15034] = 8'hd2 ;
            rom[15035] = 8'he8 ;
            rom[15036] = 8'hdd ;
            rom[15037] = 8'he4 ;
            rom[15038] = 8'hfa ;
            rom[15039] = 8'hf5 ;
            rom[15040] = 8'h2e ;
            rom[15041] = 8'h0a ;
            rom[15042] = 8'h06 ;
            rom[15043] = 8'h0d ;
            rom[15044] = 8'h11 ;
            rom[15045] = 8'hd6 ;
            rom[15046] = 8'h17 ;
            rom[15047] = 8'hea ;
            rom[15048] = 8'h01 ;
            rom[15049] = 8'hde ;
            rom[15050] = 8'hed ;
            rom[15051] = 8'hec ;
            rom[15052] = 8'h1b ;
            rom[15053] = 8'hf9 ;
            rom[15054] = 8'he9 ;
            rom[15055] = 8'h0c ;
            rom[15056] = 8'h08 ;
            rom[15057] = 8'h09 ;
            rom[15058] = 8'h1a ;
            rom[15059] = 8'h0f ;
            rom[15060] = 8'h0d ;
            rom[15061] = 8'h12 ;
            rom[15062] = 8'hfc ;
            rom[15063] = 8'h25 ;
            rom[15064] = 8'he6 ;
            rom[15065] = 8'hf4 ;
            rom[15066] = 8'hfc ;
            rom[15067] = 8'h1b ;
            rom[15068] = 8'h02 ;
            rom[15069] = 8'h1d ;
            rom[15070] = 8'hed ;
            rom[15071] = 8'hfd ;
            rom[15072] = 8'h12 ;
            rom[15073] = 8'h0c ;
            rom[15074] = 8'he3 ;
            rom[15075] = 8'h1a ;
            rom[15076] = 8'hde ;
            rom[15077] = 8'h26 ;
            rom[15078] = 8'hfa ;
            rom[15079] = 8'heb ;
            rom[15080] = 8'hf3 ;
            rom[15081] = 8'hfc ;
            rom[15082] = 8'h17 ;
            rom[15083] = 8'hfd ;
            rom[15084] = 8'h03 ;
            rom[15085] = 8'hf5 ;
            rom[15086] = 8'hde ;
            rom[15087] = 8'h14 ;
            rom[15088] = 8'hff ;
            rom[15089] = 8'hf2 ;
            rom[15090] = 8'he5 ;
            rom[15091] = 8'h1b ;
            rom[15092] = 8'hf1 ;
            rom[15093] = 8'hfa ;
            rom[15094] = 8'hf2 ;
            rom[15095] = 8'hf3 ;
            rom[15096] = 8'hee ;
            rom[15097] = 8'he9 ;
            rom[15098] = 8'hba ;
            rom[15099] = 8'hd4 ;
            rom[15100] = 8'hfb ;
            rom[15101] = 8'h09 ;
            rom[15102] = 8'hfc ;
            rom[15103] = 8'hf3 ;
            rom[15104] = 8'hf1 ;
            rom[15105] = 8'hda ;
            rom[15106] = 8'h0c ;
            rom[15107] = 8'hf7 ;
            rom[15108] = 8'he5 ;
            rom[15109] = 8'h22 ;
            rom[15110] = 8'hd3 ;
            rom[15111] = 8'hce ;
            rom[15112] = 8'h06 ;
            rom[15113] = 8'hd6 ;
            rom[15114] = 8'he4 ;
            rom[15115] = 8'heb ;
            rom[15116] = 8'h01 ;
            rom[15117] = 8'h10 ;
            rom[15118] = 8'h17 ;
            rom[15119] = 8'hed ;
            rom[15120] = 8'hf7 ;
            rom[15121] = 8'h29 ;
            rom[15122] = 8'h20 ;
            rom[15123] = 8'h03 ;
            rom[15124] = 8'he0 ;
            rom[15125] = 8'hf0 ;
            rom[15126] = 8'h12 ;
            rom[15127] = 8'h0a ;
            rom[15128] = 8'hed ;
            rom[15129] = 8'he9 ;
            rom[15130] = 8'h0e ;
            rom[15131] = 8'hed ;
            rom[15132] = 8'hef ;
            rom[15133] = 8'h0a ;
            rom[15134] = 8'h0a ;
            rom[15135] = 8'h04 ;
            rom[15136] = 8'he0 ;
            rom[15137] = 8'h09 ;
            rom[15138] = 8'hc9 ;
            rom[15139] = 8'hf7 ;
            rom[15140] = 8'hda ;
            rom[15141] = 8'hce ;
            rom[15142] = 8'h0c ;
            rom[15143] = 8'hf7 ;
            rom[15144] = 8'h03 ;
            rom[15145] = 8'h19 ;
            rom[15146] = 8'h09 ;
            rom[15147] = 8'h3b ;
            rom[15148] = 8'hd9 ;
            rom[15149] = 8'hef ;
            rom[15150] = 8'hea ;
            rom[15151] = 8'hf7 ;
            rom[15152] = 8'hf8 ;
            rom[15153] = 8'hcf ;
            rom[15154] = 8'hf3 ;
            rom[15155] = 8'h07 ;
            rom[15156] = 8'h0a ;
            rom[15157] = 8'hf5 ;
            rom[15158] = 8'h0f ;
            rom[15159] = 8'h1a ;
            rom[15160] = 8'hf4 ;
            rom[15161] = 8'h04 ;
            rom[15162] = 8'h1c ;
            rom[15163] = 8'hec ;
            rom[15164] = 8'h07 ;
            rom[15165] = 8'hde ;
            rom[15166] = 8'hea ;
            rom[15167] = 8'hfe ;
            rom[15168] = 8'h03 ;
            rom[15169] = 8'hfb ;
            rom[15170] = 8'hf0 ;
            rom[15171] = 8'hf9 ;
            rom[15172] = 8'h08 ;
            rom[15173] = 8'hf9 ;
            rom[15174] = 8'hf8 ;
            rom[15175] = 8'hfb ;
            rom[15176] = 8'hf7 ;
            rom[15177] = 8'he8 ;
            rom[15178] = 8'h04 ;
            rom[15179] = 8'hf4 ;
            rom[15180] = 8'h11 ;
            rom[15181] = 8'h03 ;
            rom[15182] = 8'hf8 ;
            rom[15183] = 8'h00 ;
            rom[15184] = 8'h07 ;
            rom[15185] = 8'hf6 ;
            rom[15186] = 8'h20 ;
            rom[15187] = 8'hd8 ;
            rom[15188] = 8'hf6 ;
            rom[15189] = 8'hf1 ;
            rom[15190] = 8'h03 ;
            rom[15191] = 8'h21 ;
            rom[15192] = 8'h0d ;
            rom[15193] = 8'h02 ;
            rom[15194] = 8'hf8 ;
            rom[15195] = 8'he1 ;
            rom[15196] = 8'hef ;
            rom[15197] = 8'he1 ;
            rom[15198] = 8'hf8 ;
            rom[15199] = 8'hfb ;
            rom[15200] = 8'hf0 ;
            rom[15201] = 8'h1a ;
            rom[15202] = 8'h0f ;
            rom[15203] = 8'he4 ;
            rom[15204] = 8'he1 ;
            rom[15205] = 8'hd2 ;
            rom[15206] = 8'h06 ;
            rom[15207] = 8'h0c ;
            rom[15208] = 8'hf0 ;
            rom[15209] = 8'h1f ;
            rom[15210] = 8'hdc ;
            rom[15211] = 8'h14 ;
            rom[15212] = 8'h1b ;
            rom[15213] = 8'hf9 ;
            rom[15214] = 8'he8 ;
            rom[15215] = 8'hf8 ;
            rom[15216] = 8'h17 ;
            rom[15217] = 8'hf7 ;
            rom[15218] = 8'h11 ;
            rom[15219] = 8'h07 ;
            rom[15220] = 8'h00 ;
            rom[15221] = 8'he2 ;
            rom[15222] = 8'hf0 ;
            rom[15223] = 8'h1f ;
            rom[15224] = 8'h03 ;
            rom[15225] = 8'h2a ;
            rom[15226] = 8'hf0 ;
            rom[15227] = 8'hf8 ;
            rom[15228] = 8'hd4 ;
            rom[15229] = 8'h0d ;
            rom[15230] = 8'h01 ;
            rom[15231] = 8'hc3 ;
            rom[15232] = 8'hf1 ;
            rom[15233] = 8'he3 ;
            rom[15234] = 8'h0c ;
            rom[15235] = 8'h15 ;
            rom[15236] = 8'h2a ;
            rom[15237] = 8'hc9 ;
            rom[15238] = 8'hf3 ;
            rom[15239] = 8'hed ;
            rom[15240] = 8'h1a ;
            rom[15241] = 8'h00 ;
            rom[15242] = 8'heb ;
            rom[15243] = 8'hff ;
            rom[15244] = 8'hcd ;
            rom[15245] = 8'hf4 ;
            rom[15246] = 8'he8 ;
            rom[15247] = 8'he6 ;
            rom[15248] = 8'hf6 ;
            rom[15249] = 8'h0a ;
            rom[15250] = 8'h20 ;
            rom[15251] = 8'h00 ;
            rom[15252] = 8'h04 ;
            rom[15253] = 8'h05 ;
            rom[15254] = 8'hf4 ;
            rom[15255] = 8'he6 ;
            rom[15256] = 8'hdf ;
            rom[15257] = 8'h1e ;
            rom[15258] = 8'h07 ;
            rom[15259] = 8'hf7 ;
            rom[15260] = 8'hfe ;
            rom[15261] = 8'h37 ;
            rom[15262] = 8'hf7 ;
            rom[15263] = 8'h17 ;
            rom[15264] = 8'h10 ;
            rom[15265] = 8'h0f ;
            rom[15266] = 8'hea ;
            rom[15267] = 8'he9 ;
            rom[15268] = 8'hd3 ;
            rom[15269] = 8'h00 ;
            rom[15270] = 8'hf9 ;
            rom[15271] = 8'h18 ;
            rom[15272] = 8'h32 ;
            rom[15273] = 8'h0c ;
            rom[15274] = 8'hf5 ;
            rom[15275] = 8'he1 ;
            rom[15276] = 8'h09 ;
            rom[15277] = 8'hfa ;
            rom[15278] = 8'hfa ;
            rom[15279] = 8'h00 ;
            rom[15280] = 8'hdf ;
            rom[15281] = 8'h00 ;
            rom[15282] = 8'h1f ;
            rom[15283] = 8'hf7 ;
            rom[15284] = 8'he5 ;
            rom[15285] = 8'he5 ;
            rom[15286] = 8'hc7 ;
            rom[15287] = 8'hf1 ;
            rom[15288] = 8'hee ;
            rom[15289] = 8'hfd ;
            rom[15290] = 8'hfd ;
            rom[15291] = 8'hd0 ;
            rom[15292] = 8'h11 ;
            rom[15293] = 8'h15 ;
            rom[15294] = 8'h1a ;
            rom[15295] = 8'he1 ;
            rom[15296] = 8'h10 ;
            rom[15297] = 8'hf1 ;
            rom[15298] = 8'h15 ;
            rom[15299] = 8'hda ;
            rom[15300] = 8'h14 ;
            rom[15301] = 8'hd9 ;
            rom[15302] = 8'hc5 ;
            rom[15303] = 8'hfd ;
            rom[15304] = 8'he4 ;
            rom[15305] = 8'h18 ;
            rom[15306] = 8'h37 ;
            rom[15307] = 8'h05 ;
            rom[15308] = 8'hf6 ;
            rom[15309] = 8'hfd ;
            rom[15310] = 8'h0b ;
            rom[15311] = 8'h15 ;
            rom[15312] = 8'hba ;
            rom[15313] = 8'h08 ;
            rom[15314] = 8'he6 ;
            rom[15315] = 8'he2 ;
            rom[15316] = 8'h05 ;
            rom[15317] = 8'h19 ;
            rom[15318] = 8'h11 ;
            rom[15319] = 8'hfd ;
            rom[15320] = 8'hf8 ;
            rom[15321] = 8'h10 ;
            rom[15322] = 8'h01 ;
            rom[15323] = 8'hf2 ;
            rom[15324] = 8'hd5 ;
            rom[15325] = 8'hfa ;
            rom[15326] = 8'h1e ;
            rom[15327] = 8'h0c ;
            rom[15328] = 8'h0d ;
            rom[15329] = 8'hf4 ;
            rom[15330] = 8'hfb ;
            rom[15331] = 8'hde ;
            rom[15332] = 8'hed ;
            rom[15333] = 8'hdd ;
            rom[15334] = 8'hca ;
            rom[15335] = 8'hc2 ;
            rom[15336] = 8'he5 ;
            rom[15337] = 8'he3 ;
            rom[15338] = 8'he9 ;
            rom[15339] = 8'h0b ;
            rom[15340] = 8'hdb ;
            rom[15341] = 8'hc9 ;
            rom[15342] = 8'hfc ;
            rom[15343] = 8'h08 ;
            rom[15344] = 8'he2 ;
            rom[15345] = 8'hfb ;
            rom[15346] = 8'h18 ;
            rom[15347] = 8'h29 ;
            rom[15348] = 8'h09 ;
            rom[15349] = 8'hfe ;
            rom[15350] = 8'h0b ;
            rom[15351] = 8'he6 ;
            rom[15352] = 8'hef ;
            rom[15353] = 8'hf4 ;
            rom[15354] = 8'hd5 ;
            rom[15355] = 8'h10 ;
            rom[15356] = 8'h10 ;
            rom[15357] = 8'hfa ;
            rom[15358] = 8'hcb ;
            rom[15359] = 8'h05 ;
            rom[15360] = 8'hf3 ;
            rom[15361] = 8'hf5 ;
            rom[15362] = 8'hf4 ;
            rom[15363] = 8'h0a ;
            rom[15364] = 8'hf4 ;
            rom[15365] = 8'hdf ;
            rom[15366] = 8'hfc ;
            rom[15367] = 8'hfc ;
            rom[15368] = 8'hfd ;
            rom[15369] = 8'hdc ;
            rom[15370] = 8'hf3 ;
            rom[15371] = 8'hfc ;
            rom[15372] = 8'h28 ;
            rom[15373] = 8'hf9 ;
            rom[15374] = 8'h0c ;
            rom[15375] = 8'hd7 ;
            rom[15376] = 8'heb ;
            rom[15377] = 8'hc2 ;
            rom[15378] = 8'hea ;
            rom[15379] = 8'h16 ;
            rom[15380] = 8'hfb ;
            rom[15381] = 8'hf4 ;
            rom[15382] = 8'he2 ;
            rom[15383] = 8'hc4 ;
            rom[15384] = 8'hea ;
            rom[15385] = 8'hf9 ;
            rom[15386] = 8'hff ;
            rom[15387] = 8'h0c ;
            rom[15388] = 8'h12 ;
            rom[15389] = 8'h08 ;
            rom[15390] = 8'hfb ;
            rom[15391] = 8'h03 ;
            rom[15392] = 8'hff ;
            rom[15393] = 8'he8 ;
            rom[15394] = 8'hfd ;
            rom[15395] = 8'hc6 ;
            rom[15396] = 8'he7 ;
            rom[15397] = 8'hf3 ;
            rom[15398] = 8'h0b ;
            rom[15399] = 8'he5 ;
            rom[15400] = 8'h05 ;
            rom[15401] = 8'he5 ;
            rom[15402] = 8'h13 ;
            rom[15403] = 8'he5 ;
            rom[15404] = 8'h04 ;
            rom[15405] = 8'h0b ;
            rom[15406] = 8'hf1 ;
            rom[15407] = 8'hfa ;
            rom[15408] = 8'h0d ;
            rom[15409] = 8'h01 ;
            rom[15410] = 8'he4 ;
            rom[15411] = 8'h01 ;
            rom[15412] = 8'hfc ;
            rom[15413] = 8'h0d ;
            rom[15414] = 8'hf4 ;
            rom[15415] = 8'he6 ;
            rom[15416] = 8'he6 ;
            rom[15417] = 8'hef ;
            rom[15418] = 8'h19 ;
            rom[15419] = 8'h1f ;
            rom[15420] = 8'h0b ;
            rom[15421] = 8'h00 ;
            rom[15422] = 8'hdd ;
            rom[15423] = 8'h01 ;
            rom[15424] = 8'h05 ;
            rom[15425] = 8'h1a ;
            rom[15426] = 8'h18 ;
            rom[15427] = 8'hf6 ;
            rom[15428] = 8'heb ;
            rom[15429] = 8'hfc ;
            rom[15430] = 8'h12 ;
            rom[15431] = 8'hf7 ;
            rom[15432] = 8'h05 ;
            rom[15433] = 8'hc6 ;
            rom[15434] = 8'hea ;
            rom[15435] = 8'h1d ;
            rom[15436] = 8'hde ;
            rom[15437] = 8'h06 ;
            rom[15438] = 8'hee ;
            rom[15439] = 8'hdf ;
            rom[15440] = 8'hf2 ;
            rom[15441] = 8'h0a ;
            rom[15442] = 8'hdc ;
            rom[15443] = 8'h0d ;
            rom[15444] = 8'h17 ;
            rom[15445] = 8'hd1 ;
            rom[15446] = 8'hf1 ;
            rom[15447] = 8'h02 ;
            rom[15448] = 8'hfe ;
            rom[15449] = 8'hd7 ;
            rom[15450] = 8'h04 ;
            rom[15451] = 8'h10 ;
            rom[15452] = 8'hce ;
            rom[15453] = 8'hf5 ;
            rom[15454] = 8'h04 ;
            rom[15455] = 8'hd2 ;
            rom[15456] = 8'he3 ;
            rom[15457] = 8'hfd ;
            rom[15458] = 8'hd7 ;
            rom[15459] = 8'h05 ;
            rom[15460] = 8'hfb ;
            rom[15461] = 8'h04 ;
            rom[15462] = 8'h0b ;
            rom[15463] = 8'hdc ;
            rom[15464] = 8'hdb ;
            rom[15465] = 8'hee ;
            rom[15466] = 8'h0a ;
            rom[15467] = 8'hfe ;
            rom[15468] = 8'hf3 ;
            rom[15469] = 8'h02 ;
            rom[15470] = 8'hfe ;
            rom[15471] = 8'h23 ;
            rom[15472] = 8'hfe ;
            rom[15473] = 8'h07 ;
            rom[15474] = 8'h11 ;
            rom[15475] = 8'h03 ;
            rom[15476] = 8'hea ;
            rom[15477] = 8'hde ;
            rom[15478] = 8'hf6 ;
            rom[15479] = 8'hce ;
            rom[15480] = 8'h29 ;
            rom[15481] = 8'he0 ;
            rom[15482] = 8'h06 ;
            rom[15483] = 8'h12 ;
            rom[15484] = 8'hf6 ;
            rom[15485] = 8'hdb ;
            rom[15486] = 8'he3 ;
            rom[15487] = 8'hdc ;
            rom[15488] = 8'hee ;
            rom[15489] = 8'heb ;
            rom[15490] = 8'h0b ;
            rom[15491] = 8'hf4 ;
            rom[15492] = 8'h19 ;
            rom[15493] = 8'hf9 ;
            rom[15494] = 8'h10 ;
            rom[15495] = 8'he3 ;
            rom[15496] = 8'h1d ;
            rom[15497] = 8'hef ;
            rom[15498] = 8'hfd ;
            rom[15499] = 8'he0 ;
            rom[15500] = 8'hdd ;
            rom[15501] = 8'he8 ;
            rom[15502] = 8'h12 ;
            rom[15503] = 8'h06 ;
            rom[15504] = 8'h10 ;
            rom[15505] = 8'h05 ;
            rom[15506] = 8'h04 ;
            rom[15507] = 8'h09 ;
            rom[15508] = 8'hf3 ;
            rom[15509] = 8'hd5 ;
            rom[15510] = 8'hd2 ;
            rom[15511] = 8'h09 ;
            rom[15512] = 8'hfe ;
            rom[15513] = 8'hee ;
            rom[15514] = 8'hfd ;
            rom[15515] = 8'hf2 ;
            rom[15516] = 8'hef ;
            rom[15517] = 8'h10 ;
            rom[15518] = 8'he8 ;
            rom[15519] = 8'h05 ;
            rom[15520] = 8'hb7 ;
            rom[15521] = 8'he0 ;
            rom[15522] = 8'hfc ;
            rom[15523] = 8'h08 ;
            rom[15524] = 8'heb ;
            rom[15525] = 8'hea ;
            rom[15526] = 8'hd8 ;
            rom[15527] = 8'hfa ;
            rom[15528] = 8'he8 ;
            rom[15529] = 8'hff ;
            rom[15530] = 8'hee ;
            rom[15531] = 8'h15 ;
            rom[15532] = 8'h0e ;
            rom[15533] = 8'h03 ;
            rom[15534] = 8'h21 ;
            rom[15535] = 8'hf0 ;
            rom[15536] = 8'hda ;
            rom[15537] = 8'hd8 ;
            rom[15538] = 8'hdf ;
            rom[15539] = 8'h0f ;
            rom[15540] = 8'h19 ;
            rom[15541] = 8'he5 ;
            rom[15542] = 8'hf6 ;
            rom[15543] = 8'hfa ;
            rom[15544] = 8'h27 ;
            rom[15545] = 8'h1e ;
            rom[15546] = 8'h0e ;
            rom[15547] = 8'hdd ;
            rom[15548] = 8'hfb ;
            rom[15549] = 8'hce ;
            rom[15550] = 8'h28 ;
            rom[15551] = 8'h0f ;
            rom[15552] = 8'he8 ;
            rom[15553] = 8'h25 ;
            rom[15554] = 8'hea ;
            rom[15555] = 8'h1d ;
            rom[15556] = 8'hea ;
            rom[15557] = 8'h02 ;
            rom[15558] = 8'hcd ;
            rom[15559] = 8'hfc ;
            rom[15560] = 8'h03 ;
            rom[15561] = 8'h11 ;
            rom[15562] = 8'heb ;
            rom[15563] = 8'he6 ;
            rom[15564] = 8'h2d ;
            rom[15565] = 8'h04 ;
            rom[15566] = 8'h2b ;
            rom[15567] = 8'hf7 ;
            rom[15568] = 8'h0a ;
            rom[15569] = 8'hf5 ;
            rom[15570] = 8'h1e ;
            rom[15571] = 8'h09 ;
            rom[15572] = 8'hda ;
            rom[15573] = 8'h15 ;
            rom[15574] = 8'he9 ;
            rom[15575] = 8'hed ;
            rom[15576] = 8'h19 ;
            rom[15577] = 8'hfe ;
            rom[15578] = 8'hf0 ;
            rom[15579] = 8'hf1 ;
            rom[15580] = 8'heb ;
            rom[15581] = 8'hfc ;
            rom[15582] = 8'h02 ;
            rom[15583] = 8'h10 ;
            rom[15584] = 8'hfc ;
            rom[15585] = 8'hd4 ;
            rom[15586] = 8'h01 ;
            rom[15587] = 8'hd6 ;
            rom[15588] = 8'hf5 ;
            rom[15589] = 8'hd6 ;
            rom[15590] = 8'h0f ;
            rom[15591] = 8'h1f ;
            rom[15592] = 8'hdd ;
            rom[15593] = 8'hf8 ;
            rom[15594] = 8'hf4 ;
            rom[15595] = 8'h08 ;
            rom[15596] = 8'hf6 ;
            rom[15597] = 8'hd6 ;
            rom[15598] = 8'h08 ;
            rom[15599] = 8'hd9 ;
            rom[15600] = 8'he7 ;
            rom[15601] = 8'hf0 ;
            rom[15602] = 8'hec ;
            rom[15603] = 8'h26 ;
            rom[15604] = 8'h14 ;
            rom[15605] = 8'h0f ;
            rom[15606] = 8'h18 ;
            rom[15607] = 8'he5 ;
            rom[15608] = 8'hf9 ;
            rom[15609] = 8'h11 ;
            rom[15610] = 8'h0a ;
            rom[15611] = 8'hf8 ;
            rom[15612] = 8'h0f ;
            rom[15613] = 8'h08 ;
            rom[15614] = 8'h17 ;
            rom[15615] = 8'h0a ;
            rom[15616] = 8'hf9 ;
            rom[15617] = 8'h01 ;
            rom[15618] = 8'h07 ;
            rom[15619] = 8'h10 ;
            rom[15620] = 8'hf5 ;
            rom[15621] = 8'hfb ;
            rom[15622] = 8'h14 ;
            rom[15623] = 8'hdc ;
            rom[15624] = 8'he8 ;
            rom[15625] = 8'h22 ;
            rom[15626] = 8'hff ;
            rom[15627] = 8'hd4 ;
            rom[15628] = 8'hdf ;
            rom[15629] = 8'h1e ;
            rom[15630] = 8'hf9 ;
            rom[15631] = 8'hda ;
            rom[15632] = 8'hd8 ;
            rom[15633] = 8'h07 ;
            rom[15634] = 8'h0b ;
            rom[15635] = 8'hfc ;
            rom[15636] = 8'hcc ;
            rom[15637] = 8'hd5 ;
            rom[15638] = 8'h3b ;
            rom[15639] = 8'h05 ;
            rom[15640] = 8'h14 ;
            rom[15641] = 8'h16 ;
            rom[15642] = 8'he7 ;
            rom[15643] = 8'h01 ;
            rom[15644] = 8'h08 ;
            rom[15645] = 8'h24 ;
            rom[15646] = 8'hec ;
            rom[15647] = 8'h04 ;
            rom[15648] = 8'he6 ;
            rom[15649] = 8'heb ;
            rom[15650] = 8'h0c ;
            rom[15651] = 8'hec ;
            rom[15652] = 8'h0c ;
            rom[15653] = 8'he5 ;
            rom[15654] = 8'h03 ;
            rom[15655] = 8'hfd ;
            rom[15656] = 8'hdb ;
            rom[15657] = 8'hdf ;
            rom[15658] = 8'he3 ;
            rom[15659] = 8'h14 ;
            rom[15660] = 8'h12 ;
            rom[15661] = 8'hd3 ;
            rom[15662] = 8'h00 ;
            rom[15663] = 8'hf7 ;
            rom[15664] = 8'h0c ;
            rom[15665] = 8'h14 ;
            rom[15666] = 8'hc4 ;
            rom[15667] = 8'hdb ;
            rom[15668] = 8'h09 ;
            rom[15669] = 8'he0 ;
            rom[15670] = 8'hfe ;
            rom[15671] = 8'h0c ;
            rom[15672] = 8'h23 ;
            rom[15673] = 8'h13 ;
            rom[15674] = 8'hf2 ;
            rom[15675] = 8'hfb ;
            rom[15676] = 8'h09 ;
            rom[15677] = 8'h03 ;
            rom[15678] = 8'h03 ;
            rom[15679] = 8'h02 ;
            rom[15680] = 8'h0a ;
            rom[15681] = 8'h00 ;
            rom[15682] = 8'h01 ;
            rom[15683] = 8'hb7 ;
            rom[15684] = 8'h1c ;
            rom[15685] = 8'hf2 ;
            rom[15686] = 8'hb8 ;
            rom[15687] = 8'h03 ;
            rom[15688] = 8'hfb ;
            rom[15689] = 8'hfe ;
            rom[15690] = 8'hf5 ;
            rom[15691] = 8'hdf ;
            rom[15692] = 8'he8 ;
            rom[15693] = 8'he0 ;
            rom[15694] = 8'hf2 ;
            rom[15695] = 8'h1d ;
            rom[15696] = 8'h0e ;
            rom[15697] = 8'h11 ;
            rom[15698] = 8'h19 ;
            rom[15699] = 8'hf8 ;
            rom[15700] = 8'hf3 ;
            rom[15701] = 8'h15 ;
            rom[15702] = 8'he0 ;
            rom[15703] = 8'hed ;
            rom[15704] = 8'he0 ;
            rom[15705] = 8'hd1 ;
            rom[15706] = 8'hc4 ;
            rom[15707] = 8'h25 ;
            rom[15708] = 8'hfa ;
            rom[15709] = 8'hf4 ;
            rom[15710] = 8'hed ;
            rom[15711] = 8'hfb ;
            rom[15712] = 8'h08 ;
            rom[15713] = 8'hed ;
            rom[15714] = 8'h08 ;
            rom[15715] = 8'h1a ;
            rom[15716] = 8'h0b ;
            rom[15717] = 8'h17 ;
            rom[15718] = 8'h0b ;
            rom[15719] = 8'hf3 ;
            rom[15720] = 8'hbf ;
            rom[15721] = 8'h00 ;
            rom[15722] = 8'h18 ;
            rom[15723] = 8'h25 ;
            rom[15724] = 8'hff ;
            rom[15725] = 8'hf2 ;
            rom[15726] = 8'h0f ;
            rom[15727] = 8'he5 ;
            rom[15728] = 8'hdd ;
            rom[15729] = 8'hf3 ;
            rom[15730] = 8'h0c ;
            rom[15731] = 8'h0b ;
            rom[15732] = 8'h07 ;
            rom[15733] = 8'hfe ;
            rom[15734] = 8'hf5 ;
            rom[15735] = 8'h08 ;
            rom[15736] = 8'hdc ;
            rom[15737] = 8'h03 ;
            rom[15738] = 8'hf4 ;
            rom[15739] = 8'h0e ;
            rom[15740] = 8'hda ;
            rom[15741] = 8'h1b ;
            rom[15742] = 8'h08 ;
            rom[15743] = 8'h14 ;
            rom[15744] = 8'hf0 ;
            rom[15745] = 8'hf6 ;
            rom[15746] = 8'hf4 ;
            rom[15747] = 8'h09 ;
            rom[15748] = 8'h24 ;
            rom[15749] = 8'hbd ;
            rom[15750] = 8'hf0 ;
            rom[15751] = 8'hd9 ;
            rom[15752] = 8'he2 ;
            rom[15753] = 8'hf6 ;
            rom[15754] = 8'he0 ;
            rom[15755] = 8'hf4 ;
            rom[15756] = 8'hcb ;
            rom[15757] = 8'hf0 ;
            rom[15758] = 8'he5 ;
            rom[15759] = 8'hff ;
            rom[15760] = 8'hef ;
            rom[15761] = 8'h1a ;
            rom[15762] = 8'h04 ;
            rom[15763] = 8'hcf ;
            rom[15764] = 8'h07 ;
            rom[15765] = 8'h0c ;
            rom[15766] = 8'hfd ;
            rom[15767] = 8'h1d ;
            rom[15768] = 8'he3 ;
            rom[15769] = 8'hf1 ;
            rom[15770] = 8'h0b ;
            rom[15771] = 8'hfe ;
            rom[15772] = 8'hf2 ;
            rom[15773] = 8'h18 ;
            rom[15774] = 8'hd7 ;
            rom[15775] = 8'h0c ;
            rom[15776] = 8'h0f ;
            rom[15777] = 8'he7 ;
            rom[15778] = 8'h0c ;
            rom[15779] = 8'hbe ;
            rom[15780] = 8'hdd ;
            rom[15781] = 8'hcb ;
            rom[15782] = 8'hf2 ;
            rom[15783] = 8'h05 ;
            rom[15784] = 8'h24 ;
            rom[15785] = 8'hef ;
            rom[15786] = 8'hf9 ;
            rom[15787] = 8'h1f ;
            rom[15788] = 8'hf1 ;
            rom[15789] = 8'hcb ;
            rom[15790] = 8'h06 ;
            rom[15791] = 8'h08 ;
            rom[15792] = 8'h04 ;
            rom[15793] = 8'hfb ;
            rom[15794] = 8'h01 ;
            rom[15795] = 8'h09 ;
            rom[15796] = 8'h16 ;
            rom[15797] = 8'h0a ;
            rom[15798] = 8'h0c ;
            rom[15799] = 8'he2 ;
            rom[15800] = 8'h1f ;
            rom[15801] = 8'hf0 ;
            rom[15802] = 8'h09 ;
            rom[15803] = 8'h0a ;
            rom[15804] = 8'hf2 ;
            rom[15805] = 8'h02 ;
            rom[15806] = 8'h09 ;
            rom[15807] = 8'hec ;
            rom[15808] = 8'hf4 ;
            rom[15809] = 8'h08 ;
            rom[15810] = 8'hc5 ;
            rom[15811] = 8'h08 ;
            rom[15812] = 8'hf9 ;
            rom[15813] = 8'h10 ;
            rom[15814] = 8'he4 ;
            rom[15815] = 8'hee ;
            rom[15816] = 8'h0a ;
            rom[15817] = 8'he9 ;
            rom[15818] = 8'h09 ;
            rom[15819] = 8'he2 ;
            rom[15820] = 8'hdd ;
            rom[15821] = 8'hd0 ;
            rom[15822] = 8'he1 ;
            rom[15823] = 8'h0c ;
            rom[15824] = 8'hd7 ;
            rom[15825] = 8'hf0 ;
            rom[15826] = 8'h1e ;
            rom[15827] = 8'h05 ;
            rom[15828] = 8'hed ;
            rom[15829] = 8'hf4 ;
            rom[15830] = 8'hec ;
            rom[15831] = 8'hf8 ;
            rom[15832] = 8'hff ;
            rom[15833] = 8'h18 ;
            rom[15834] = 8'h20 ;
            rom[15835] = 8'h10 ;
            rom[15836] = 8'hf9 ;
            rom[15837] = 8'h09 ;
            rom[15838] = 8'h0a ;
            rom[15839] = 8'h08 ;
            rom[15840] = 8'h04 ;
            rom[15841] = 8'hf2 ;
            rom[15842] = 8'h06 ;
            rom[15843] = 8'hd7 ;
            rom[15844] = 8'h09 ;
            rom[15845] = 8'hdb ;
            rom[15846] = 8'h10 ;
            rom[15847] = 8'h17 ;
            rom[15848] = 8'hef ;
            rom[15849] = 8'hf7 ;
            rom[15850] = 8'he7 ;
            rom[15851] = 8'h25 ;
            rom[15852] = 8'hd5 ;
            rom[15853] = 8'he2 ;
            rom[15854] = 8'hc6 ;
            rom[15855] = 8'h22 ;
            rom[15856] = 8'hf2 ;
            rom[15857] = 8'h0a ;
            rom[15858] = 8'hd3 ;
            rom[15859] = 8'h10 ;
            rom[15860] = 8'h18 ;
            rom[15861] = 8'hf2 ;
            rom[15862] = 8'h19 ;
            rom[15863] = 8'heb ;
            rom[15864] = 8'h11 ;
            rom[15865] = 8'h28 ;
            rom[15866] = 8'hf8 ;
            rom[15867] = 8'hfd ;
            rom[15868] = 8'h1f ;
            rom[15869] = 8'h16 ;
            rom[15870] = 8'hff ;
            rom[15871] = 8'hf4 ;
            rom[15872] = 8'hf5 ;
            rom[15873] = 8'hf0 ;
            rom[15874] = 8'hdb ;
            rom[15875] = 8'h25 ;
            rom[15876] = 8'h0a ;
            rom[15877] = 8'hdf ;
            rom[15878] = 8'hf7 ;
            rom[15879] = 8'hbf ;
            rom[15880] = 8'hf0 ;
            rom[15881] = 8'h02 ;
            rom[15882] = 8'h02 ;
            rom[15883] = 8'hdb ;
            rom[15884] = 8'he4 ;
            rom[15885] = 8'hf1 ;
            rom[15886] = 8'hfa ;
            rom[15887] = 8'hd2 ;
            rom[15888] = 8'hde ;
            rom[15889] = 8'h22 ;
            rom[15890] = 8'h0c ;
            rom[15891] = 8'hf1 ;
            rom[15892] = 8'h0c ;
            rom[15893] = 8'he9 ;
            rom[15894] = 8'he8 ;
            rom[15895] = 8'h06 ;
            rom[15896] = 8'h11 ;
            rom[15897] = 8'hfe ;
            rom[15898] = 8'h09 ;
            rom[15899] = 8'hf5 ;
            rom[15900] = 8'hc5 ;
            rom[15901] = 8'h22 ;
            rom[15902] = 8'hff ;
            rom[15903] = 8'h06 ;
            rom[15904] = 8'hf3 ;
            rom[15905] = 8'hf1 ;
            rom[15906] = 8'heb ;
            rom[15907] = 8'hea ;
            rom[15908] = 8'hd6 ;
            rom[15909] = 8'hea ;
            rom[15910] = 8'hed ;
            rom[15911] = 8'h12 ;
            rom[15912] = 8'hca ;
            rom[15913] = 8'hb8 ;
            rom[15914] = 8'hec ;
            rom[15915] = 8'hfc ;
            rom[15916] = 8'hff ;
            rom[15917] = 8'hf2 ;
            rom[15918] = 8'h04 ;
            rom[15919] = 8'hfa ;
            rom[15920] = 8'hd3 ;
            rom[15921] = 8'h04 ;
            rom[15922] = 8'h00 ;
            rom[15923] = 8'hec ;
            rom[15924] = 8'h0c ;
            rom[15925] = 8'he3 ;
            rom[15926] = 8'hf5 ;
            rom[15927] = 8'h0c ;
            rom[15928] = 8'h11 ;
            rom[15929] = 8'hfb ;
            rom[15930] = 8'h10 ;
            rom[15931] = 8'hb0 ;
            rom[15932] = 8'h05 ;
            rom[15933] = 8'hc8 ;
            rom[15934] = 8'h04 ;
            rom[15935] = 8'hd1 ;
            rom[15936] = 8'hda ;
            rom[15937] = 8'hfe ;
            rom[15938] = 8'h05 ;
            rom[15939] = 8'h03 ;
            rom[15940] = 8'h09 ;
            rom[15941] = 8'hf1 ;
            rom[15942] = 8'h04 ;
            rom[15943] = 8'he3 ;
            rom[15944] = 8'he3 ;
            rom[15945] = 8'hca ;
            rom[15946] = 8'h0a ;
            rom[15947] = 8'h28 ;
            rom[15948] = 8'h0b ;
            rom[15949] = 8'h0a ;
            rom[15950] = 8'h13 ;
            rom[15951] = 8'h03 ;
            rom[15952] = 8'hd8 ;
            rom[15953] = 8'he4 ;
            rom[15954] = 8'hf0 ;
            rom[15955] = 8'hd6 ;
            rom[15956] = 8'hd9 ;
            rom[15957] = 8'hf6 ;
            rom[15958] = 8'he4 ;
            rom[15959] = 8'hf5 ;
            rom[15960] = 8'h02 ;
            rom[15961] = 8'h0c ;
            rom[15962] = 8'heb ;
            rom[15963] = 8'h16 ;
            rom[15964] = 8'h15 ;
            rom[15965] = 8'h02 ;
            rom[15966] = 8'h03 ;
            rom[15967] = 8'he6 ;
            rom[15968] = 8'hef ;
            rom[15969] = 8'hf0 ;
            rom[15970] = 8'h07 ;
            rom[15971] = 8'he0 ;
            rom[15972] = 8'hea ;
            rom[15973] = 8'hf5 ;
            rom[15974] = 8'hfd ;
            rom[15975] = 8'hf6 ;
            rom[15976] = 8'hff ;
            rom[15977] = 8'hf6 ;
            rom[15978] = 8'heb ;
            rom[15979] = 8'hff ;
            rom[15980] = 8'hd8 ;
            rom[15981] = 8'h11 ;
            rom[15982] = 8'hfd ;
            rom[15983] = 8'h08 ;
            rom[15984] = 8'hff ;
            rom[15985] = 8'h10 ;
            rom[15986] = 8'h1d ;
            rom[15987] = 8'h00 ;
            rom[15988] = 8'h13 ;
            rom[15989] = 8'h00 ;
            rom[15990] = 8'h2a ;
            rom[15991] = 8'h1a ;
            rom[15992] = 8'he8 ;
            rom[15993] = 8'h1d ;
            rom[15994] = 8'h02 ;
            rom[15995] = 8'hf3 ;
            rom[15996] = 8'hf9 ;
            rom[15997] = 8'hfc ;
            rom[15998] = 8'hea ;
            rom[15999] = 8'he6 ;
            rom[16000] = 8'he8 ;
            rom[16001] = 8'hfa ;
            rom[16002] = 8'hef ;
            rom[16003] = 8'hda ;
            rom[16004] = 8'hfd ;
            rom[16005] = 8'hee ;
            rom[16006] = 8'h09 ;
            rom[16007] = 8'hf7 ;
            rom[16008] = 8'hd2 ;
            rom[16009] = 8'hfa ;
            rom[16010] = 8'h06 ;
            rom[16011] = 8'he4 ;
            rom[16012] = 8'he7 ;
            rom[16013] = 8'hfd ;
            rom[16014] = 8'he8 ;
            rom[16015] = 8'hd3 ;
            rom[16016] = 8'h10 ;
            rom[16017] = 8'hf3 ;
            rom[16018] = 8'hee ;
            rom[16019] = 8'h05 ;
            rom[16020] = 8'he2 ;
            rom[16021] = 8'h03 ;
            rom[16022] = 8'h13 ;
            rom[16023] = 8'he8 ;
            rom[16024] = 8'hff ;
            rom[16025] = 8'h03 ;
            rom[16026] = 8'hf2 ;
            rom[16027] = 8'hcf ;
            rom[16028] = 8'he6 ;
            rom[16029] = 8'h18 ;
            rom[16030] = 8'h02 ;
            rom[16031] = 8'h17 ;
            rom[16032] = 8'h17 ;
            rom[16033] = 8'heb ;
            rom[16034] = 8'h05 ;
            rom[16035] = 8'hf7 ;
            rom[16036] = 8'h0f ;
            rom[16037] = 8'h08 ;
            rom[16038] = 8'he4 ;
            rom[16039] = 8'he7 ;
            rom[16040] = 8'hf9 ;
            rom[16041] = 8'he5 ;
            rom[16042] = 8'hdd ;
            rom[16043] = 8'h00 ;
            rom[16044] = 8'hf2 ;
            rom[16045] = 8'he4 ;
            rom[16046] = 8'hf4 ;
            rom[16047] = 8'h0c ;
            rom[16048] = 8'h05 ;
            rom[16049] = 8'hed ;
            rom[16050] = 8'hf6 ;
            rom[16051] = 8'h00 ;
            rom[16052] = 8'hc6 ;
            rom[16053] = 8'hf3 ;
            rom[16054] = 8'h0c ;
            rom[16055] = 8'hed ;
            rom[16056] = 8'hfb ;
            rom[16057] = 8'h21 ;
            rom[16058] = 8'hf4 ;
            rom[16059] = 8'hfd ;
            rom[16060] = 8'h25 ;
            rom[16061] = 8'hdd ;
            rom[16062] = 8'h00 ;
            rom[16063] = 8'h0f ;
            rom[16064] = 8'h17 ;
            rom[16065] = 8'h08 ;
            rom[16066] = 8'h15 ;
            rom[16067] = 8'hd2 ;
            rom[16068] = 8'hfa ;
            rom[16069] = 8'h0f ;
            rom[16070] = 8'hd6 ;
            rom[16071] = 8'hf9 ;
            rom[16072] = 8'hf1 ;
            rom[16073] = 8'h23 ;
            rom[16074] = 8'hc3 ;
            rom[16075] = 8'he5 ;
            rom[16076] = 8'he1 ;
            rom[16077] = 8'hb8 ;
            rom[16078] = 8'h05 ;
            rom[16079] = 8'h02 ;
            rom[16080] = 8'h0e ;
            rom[16081] = 8'h08 ;
            rom[16082] = 8'hfa ;
            rom[16083] = 8'hd5 ;
            rom[16084] = 8'hed ;
            rom[16085] = 8'hf3 ;
            rom[16086] = 8'hd3 ;
            rom[16087] = 8'h02 ;
            rom[16088] = 8'hfb ;
            rom[16089] = 8'h06 ;
            rom[16090] = 8'he2 ;
            rom[16091] = 8'he6 ;
            rom[16092] = 8'hdd ;
            rom[16093] = 8'h12 ;
            rom[16094] = 8'he2 ;
            rom[16095] = 8'hef ;
            rom[16096] = 8'hea ;
            rom[16097] = 8'hff ;
            rom[16098] = 8'hf4 ;
            rom[16099] = 8'hf0 ;
            rom[16100] = 8'hfa ;
            rom[16101] = 8'h29 ;
            rom[16102] = 8'h1b ;
            rom[16103] = 8'hd9 ;
            rom[16104] = 8'h0f ;
            rom[16105] = 8'hfe ;
            rom[16106] = 8'h0d ;
            rom[16107] = 8'hef ;
            rom[16108] = 8'he4 ;
            rom[16109] = 8'hf1 ;
            rom[16110] = 8'h2a ;
            rom[16111] = 8'heb ;
            rom[16112] = 8'hef ;
            rom[16113] = 8'hf3 ;
            rom[16114] = 8'hff ;
            rom[16115] = 8'hf6 ;
            rom[16116] = 8'h0d ;
            rom[16117] = 8'h09 ;
            rom[16118] = 8'hdb ;
            rom[16119] = 8'hff ;
            rom[16120] = 8'hf7 ;
            rom[16121] = 8'h0d ;
            rom[16122] = 8'hd6 ;
            rom[16123] = 8'hfc ;
            rom[16124] = 8'hdd ;
            rom[16125] = 8'h0d ;
            rom[16126] = 8'hf6 ;
            rom[16127] = 8'h13 ;
            rom[16128] = 8'hf0 ;
            rom[16129] = 8'hf2 ;
            rom[16130] = 8'hf3 ;
            rom[16131] = 8'h04 ;
            rom[16132] = 8'h00 ;
            rom[16133] = 8'h09 ;
            rom[16134] = 8'hf4 ;
            rom[16135] = 8'h15 ;
            rom[16136] = 8'hf2 ;
            rom[16137] = 8'h00 ;
            rom[16138] = 8'he8 ;
            rom[16139] = 8'hf2 ;
            rom[16140] = 8'hcc ;
            rom[16141] = 8'hed ;
            rom[16142] = 8'hff ;
            rom[16143] = 8'h22 ;
            rom[16144] = 8'h07 ;
            rom[16145] = 8'he9 ;
            rom[16146] = 8'hfd ;
            rom[16147] = 8'he9 ;
            rom[16148] = 8'h10 ;
            rom[16149] = 8'he5 ;
            rom[16150] = 8'hd4 ;
            rom[16151] = 8'h12 ;
            rom[16152] = 8'he8 ;
            rom[16153] = 8'h0f ;
            rom[16154] = 8'h04 ;
            rom[16155] = 8'h00 ;
            rom[16156] = 8'he4 ;
            rom[16157] = 8'h06 ;
            rom[16158] = 8'hf6 ;
            rom[16159] = 8'hc3 ;
            rom[16160] = 8'hf4 ;
            rom[16161] = 8'h10 ;
            rom[16162] = 8'h14 ;
            rom[16163] = 8'h1d ;
            rom[16164] = 8'hcd ;
            rom[16165] = 8'h07 ;
            rom[16166] = 8'h04 ;
            rom[16167] = 8'hf6 ;
            rom[16168] = 8'hdf ;
            rom[16169] = 8'he2 ;
            rom[16170] = 8'hee ;
            rom[16171] = 8'h27 ;
            rom[16172] = 8'hf6 ;
            rom[16173] = 8'hf4 ;
            rom[16174] = 8'h0f ;
            rom[16175] = 8'hf8 ;
            rom[16176] = 8'hd2 ;
            rom[16177] = 8'hd8 ;
            rom[16178] = 8'hec ;
            rom[16179] = 8'he3 ;
            rom[16180] = 8'h00 ;
            rom[16181] = 8'h00 ;
            rom[16182] = 8'hdb ;
            rom[16183] = 8'h06 ;
            rom[16184] = 8'h0c ;
            rom[16185] = 8'he9 ;
            rom[16186] = 8'hf4 ;
            rom[16187] = 8'hd1 ;
            rom[16188] = 8'hfa ;
            rom[16189] = 8'hd4 ;
            rom[16190] = 8'h0f ;
            rom[16191] = 8'hef ;
            rom[16192] = 8'hd2 ;
            rom[16193] = 8'hfc ;
            rom[16194] = 8'hef ;
            rom[16195] = 8'h1f ;
            rom[16196] = 8'hf0 ;
            rom[16197] = 8'hec ;
            rom[16198] = 8'h09 ;
            rom[16199] = 8'h00 ;
            rom[16200] = 8'hcc ;
            rom[16201] = 8'hf4 ;
            rom[16202] = 8'h00 ;
            rom[16203] = 8'h08 ;
            rom[16204] = 8'h21 ;
            rom[16205] = 8'he4 ;
            rom[16206] = 8'h04 ;
            rom[16207] = 8'h24 ;
            rom[16208] = 8'he4 ;
            rom[16209] = 8'he7 ;
            rom[16210] = 8'h12 ;
            rom[16211] = 8'hf9 ;
            rom[16212] = 8'he8 ;
            rom[16213] = 8'hf6 ;
            rom[16214] = 8'he6 ;
            rom[16215] = 8'h14 ;
            rom[16216] = 8'h20 ;
            rom[16217] = 8'h11 ;
            rom[16218] = 8'h0d ;
            rom[16219] = 8'h16 ;
            rom[16220] = 8'h01 ;
            rom[16221] = 8'h04 ;
            rom[16222] = 8'h15 ;
            rom[16223] = 8'hfe ;
            rom[16224] = 8'hfd ;
            rom[16225] = 8'hed ;
            rom[16226] = 8'hf4 ;
            rom[16227] = 8'he6 ;
            rom[16228] = 8'he1 ;
            rom[16229] = 8'hf4 ;
            rom[16230] = 8'h09 ;
            rom[16231] = 8'h17 ;
            rom[16232] = 8'hee ;
            rom[16233] = 8'hee ;
            rom[16234] = 8'h21 ;
            rom[16235] = 8'hed ;
            rom[16236] = 8'h0f ;
            rom[16237] = 8'hec ;
            rom[16238] = 8'hfa ;
            rom[16239] = 8'he4 ;
            rom[16240] = 8'h0b ;
            rom[16241] = 8'h04 ;
            rom[16242] = 8'h0e ;
            rom[16243] = 8'h15 ;
            rom[16244] = 8'h0b ;
            rom[16245] = 8'hf9 ;
            rom[16246] = 8'h22 ;
            rom[16247] = 8'hef ;
            rom[16248] = 8'hf9 ;
            rom[16249] = 8'hf3 ;
            rom[16250] = 8'h19 ;
            rom[16251] = 8'h0a ;
            rom[16252] = 8'h06 ;
            rom[16253] = 8'he9 ;
            rom[16254] = 8'h07 ;
            rom[16255] = 8'hda ;
            rom[16256] = 8'hf4 ;
            rom[16257] = 8'h13 ;
            rom[16258] = 8'hec ;
            rom[16259] = 8'hcb ;
            rom[16260] = 8'h0e ;
            rom[16261] = 8'h01 ;
            rom[16262] = 8'h28 ;
            rom[16263] = 8'h23 ;
            rom[16264] = 8'he5 ;
            rom[16265] = 8'h18 ;
            rom[16266] = 8'hde ;
            rom[16267] = 8'h00 ;
            rom[16268] = 8'h0c ;
            rom[16269] = 8'h03 ;
            rom[16270] = 8'h0c ;
            rom[16271] = 8'he8 ;
            rom[16272] = 8'h0d ;
            rom[16273] = 8'hed ;
            rom[16274] = 8'h03 ;
            rom[16275] = 8'h09 ;
            rom[16276] = 8'he3 ;
            rom[16277] = 8'hd1 ;
            rom[16278] = 8'h09 ;
            rom[16279] = 8'hdb ;
            rom[16280] = 8'he2 ;
            rom[16281] = 8'h07 ;
            rom[16282] = 8'ha7 ;
            rom[16283] = 8'hc9 ;
            rom[16284] = 8'h17 ;
            rom[16285] = 8'hbd ;
            rom[16286] = 8'hb3 ;
            rom[16287] = 8'hda ;
            rom[16288] = 8'he1 ;
            rom[16289] = 8'hee ;
            rom[16290] = 8'h05 ;
            rom[16291] = 8'h0f ;
            rom[16292] = 8'h18 ;
            rom[16293] = 8'he3 ;
            rom[16294] = 8'h06 ;
            rom[16295] = 8'h0c ;
            rom[16296] = 8'h19 ;
            rom[16297] = 8'hfd ;
            rom[16298] = 8'h05 ;
            rom[16299] = 8'hca ;
            rom[16300] = 8'hdb ;
            rom[16301] = 8'hfc ;
            rom[16302] = 8'h11 ;
            rom[16303] = 8'hc7 ;
            rom[16304] = 8'h0c ;
            rom[16305] = 8'h03 ;
            rom[16306] = 8'hf7 ;
            rom[16307] = 8'hf0 ;
            rom[16308] = 8'h03 ;
            rom[16309] = 8'h06 ;
            rom[16310] = 8'hf7 ;
            rom[16311] = 8'h10 ;
            rom[16312] = 8'hfa ;
            rom[16313] = 8'h19 ;
            rom[16314] = 8'hd8 ;
            rom[16315] = 8'hec ;
            rom[16316] = 8'h01 ;
            rom[16317] = 8'hbc ;
            rom[16318] = 8'hc1 ;
            rom[16319] = 8'h17 ;
            rom[16320] = 8'h20 ;
            rom[16321] = 8'h0b ;
            rom[16322] = 8'hf7 ;
            rom[16323] = 8'hda ;
            rom[16324] = 8'hf9 ;
            rom[16325] = 8'h01 ;
            rom[16326] = 8'hf7 ;
            rom[16327] = 8'h0f ;
            rom[16328] = 8'hef ;
            rom[16329] = 8'h02 ;
            rom[16330] = 8'hfc ;
            rom[16331] = 8'h0b ;
            rom[16332] = 8'h01 ;
            rom[16333] = 8'he7 ;
            rom[16334] = 8'heb ;
            rom[16335] = 8'h05 ;
            rom[16336] = 8'h0f ;
            rom[16337] = 8'hde ;
            rom[16338] = 8'hda ;
            rom[16339] = 8'h01 ;
            rom[16340] = 8'hf8 ;
            rom[16341] = 8'h1f ;
            rom[16342] = 8'he0 ;
            rom[16343] = 8'h15 ;
            rom[16344] = 8'he4 ;
            rom[16345] = 8'hda ;
            rom[16346] = 8'he3 ;
            rom[16347] = 8'hd4 ;
            rom[16348] = 8'hd6 ;
            rom[16349] = 8'hdb ;
            rom[16350] = 8'hc4 ;
            rom[16351] = 8'hfe ;
            rom[16352] = 8'hfe ;
            rom[16353] = 8'hd6 ;
            rom[16354] = 8'h04 ;
            rom[16355] = 8'h18 ;
            rom[16356] = 8'hf9 ;
            rom[16357] = 8'h04 ;
            rom[16358] = 8'he8 ;
            rom[16359] = 8'h20 ;
            rom[16360] = 8'hf8 ;
            rom[16361] = 8'h02 ;
            rom[16362] = 8'hfb ;
            rom[16363] = 8'hd0 ;
            rom[16364] = 8'h2a ;
            rom[16365] = 8'hf3 ;
            rom[16366] = 8'hff ;
            rom[16367] = 8'hea ;
            rom[16368] = 8'heb ;
            rom[16369] = 8'hf0 ;
            rom[16370] = 8'h0b ;
            rom[16371] = 8'hd6 ;
            rom[16372] = 8'h04 ;
            rom[16373] = 8'hef ;
            rom[16374] = 8'hfc ;
            rom[16375] = 8'h07 ;
            rom[16376] = 8'hff ;
            rom[16377] = 8'h01 ;
            rom[16378] = 8'he9 ;
            rom[16379] = 8'hf9 ;
            rom[16380] = 8'hee ;
            rom[16381] = 8'hfe ;
            rom[16382] = 8'hf9 ;
            rom[16383] = 8'h07 ;
            rom[16384] = 8'he5 ;
            rom[16385] = 8'h01 ;
            rom[16386] = 8'hf4 ;
            rom[16387] = 8'h00 ;
            rom[16388] = 8'h2a ;
            rom[16389] = 8'h16 ;
            rom[16390] = 8'h12 ;
            rom[16391] = 8'hcb ;
            rom[16392] = 8'h00 ;
            rom[16393] = 8'he2 ;
            rom[16394] = 8'h24 ;
            rom[16395] = 8'h1c ;
            rom[16396] = 8'h1c ;
            rom[16397] = 8'hec ;
            rom[16398] = 8'h00 ;
            rom[16399] = 8'h12 ;
            rom[16400] = 8'h0f ;
            rom[16401] = 8'hed ;
            rom[16402] = 8'hfa ;
            rom[16403] = 8'hdb ;
            rom[16404] = 8'h1b ;
            rom[16405] = 8'hf7 ;
            rom[16406] = 8'hf4 ;
            rom[16407] = 8'hdc ;
            rom[16408] = 8'h11 ;
            rom[16409] = 8'h02 ;
            rom[16410] = 8'hd9 ;
            rom[16411] = 8'h04 ;
            rom[16412] = 8'h05 ;
            rom[16413] = 8'h03 ;
            rom[16414] = 8'h07 ;
            rom[16415] = 8'h11 ;
            rom[16416] = 8'h01 ;
            rom[16417] = 8'hfa ;
            rom[16418] = 8'heb ;
            rom[16419] = 8'hff ;
            rom[16420] = 8'hff ;
            rom[16421] = 8'h24 ;
            rom[16422] = 8'hf6 ;
            rom[16423] = 8'h11 ;
            rom[16424] = 8'he0 ;
            rom[16425] = 8'h0c ;
            rom[16426] = 8'hf2 ;
            rom[16427] = 8'h09 ;
            rom[16428] = 8'h02 ;
            rom[16429] = 8'h34 ;
            rom[16430] = 8'h21 ;
            rom[16431] = 8'hc8 ;
            rom[16432] = 8'hf9 ;
            rom[16433] = 8'hf6 ;
            rom[16434] = 8'hbe ;
            rom[16435] = 8'hfe ;
            rom[16436] = 8'he6 ;
            rom[16437] = 8'hf9 ;
            rom[16438] = 8'hd5 ;
            rom[16439] = 8'hfd ;
            rom[16440] = 8'h06 ;
            rom[16441] = 8'h11 ;
            rom[16442] = 8'hf9 ;
            rom[16443] = 8'h0d ;
            rom[16444] = 8'h16 ;
            rom[16445] = 8'heb ;
            rom[16446] = 8'h0c ;
            rom[16447] = 8'hfd ;
            rom[16448] = 8'hf4 ;
            rom[16449] = 8'he0 ;
            rom[16450] = 8'he2 ;
            rom[16451] = 8'h2f ;
            rom[16452] = 8'he4 ;
            rom[16453] = 8'hf4 ;
            rom[16454] = 8'hd4 ;
            rom[16455] = 8'h11 ;
            rom[16456] = 8'h0b ;
            rom[16457] = 8'hf6 ;
            rom[16458] = 8'hfc ;
            rom[16459] = 8'hfd ;
            rom[16460] = 8'he6 ;
            rom[16461] = 8'haa ;
            rom[16462] = 8'h03 ;
            rom[16463] = 8'he9 ;
            rom[16464] = 8'h18 ;
            rom[16465] = 8'hfa ;
            rom[16466] = 8'h06 ;
            rom[16467] = 8'h1c ;
            rom[16468] = 8'hec ;
            rom[16469] = 8'hfc ;
            rom[16470] = 8'hfa ;
            rom[16471] = 8'h0e ;
            rom[16472] = 8'h1f ;
            rom[16473] = 8'h0c ;
            rom[16474] = 8'hfd ;
            rom[16475] = 8'hfd ;
            rom[16476] = 8'h1a ;
            rom[16477] = 8'hf7 ;
            rom[16478] = 8'h0a ;
            rom[16479] = 8'h02 ;
            rom[16480] = 8'hda ;
            rom[16481] = 8'hea ;
            rom[16482] = 8'hfd ;
            rom[16483] = 8'hc1 ;
            rom[16484] = 8'hfb ;
            rom[16485] = 8'h06 ;
            rom[16486] = 8'h2c ;
            rom[16487] = 8'hd0 ;
            rom[16488] = 8'he4 ;
            rom[16489] = 8'h29 ;
            rom[16490] = 8'hd5 ;
            rom[16491] = 8'he1 ;
            rom[16492] = 8'hf7 ;
            rom[16493] = 8'hd4 ;
            rom[16494] = 8'hfc ;
            rom[16495] = 8'h16 ;
            rom[16496] = 8'hf8 ;
            rom[16497] = 8'hea ;
            rom[16498] = 8'h2a ;
            rom[16499] = 8'h05 ;
            rom[16500] = 8'hff ;
            rom[16501] = 8'h3d ;
            rom[16502] = 8'hf3 ;
            rom[16503] = 8'hf4 ;
            rom[16504] = 8'h11 ;
            rom[16505] = 8'he0 ;
            rom[16506] = 8'hff ;
            rom[16507] = 8'he9 ;
            rom[16508] = 8'he1 ;
            rom[16509] = 8'h13 ;
            rom[16510] = 8'hfa ;
            rom[16511] = 8'he2 ;
            rom[16512] = 8'h06 ;
            rom[16513] = 8'hff ;
            rom[16514] = 8'hef ;
            rom[16515] = 8'hff ;
            rom[16516] = 8'h0c ;
            rom[16517] = 8'hd1 ;
            rom[16518] = 8'he6 ;
            rom[16519] = 8'he0 ;
            rom[16520] = 8'he6 ;
            rom[16521] = 8'h0b ;
            rom[16522] = 8'hfd ;
            rom[16523] = 8'h14 ;
            rom[16524] = 8'h04 ;
            rom[16525] = 8'h00 ;
            rom[16526] = 8'he3 ;
            rom[16527] = 8'hc3 ;
            rom[16528] = 8'hf8 ;
            rom[16529] = 8'hfa ;
            rom[16530] = 8'hdb ;
            rom[16531] = 8'hf7 ;
            rom[16532] = 8'h00 ;
            rom[16533] = 8'hdf ;
            rom[16534] = 8'hf3 ;
            rom[16535] = 8'hb3 ;
            rom[16536] = 8'hee ;
            rom[16537] = 8'h01 ;
            rom[16538] = 8'he6 ;
            rom[16539] = 8'hd4 ;
            rom[16540] = 8'hf9 ;
            rom[16541] = 8'hdb ;
            rom[16542] = 8'heb ;
            rom[16543] = 8'hf2 ;
            rom[16544] = 8'he2 ;
            rom[16545] = 8'h2b ;
            rom[16546] = 8'he2 ;
            rom[16547] = 8'h15 ;
            rom[16548] = 8'hfe ;
            rom[16549] = 8'he9 ;
            rom[16550] = 8'hfc ;
            rom[16551] = 8'hf3 ;
            rom[16552] = 8'h07 ;
            rom[16553] = 8'he3 ;
            rom[16554] = 8'he9 ;
            rom[16555] = 8'he8 ;
            rom[16556] = 8'hf1 ;
            rom[16557] = 8'he1 ;
            rom[16558] = 8'he9 ;
            rom[16559] = 8'h07 ;
            rom[16560] = 8'heb ;
            rom[16561] = 8'h0a ;
            rom[16562] = 8'h11 ;
            rom[16563] = 8'hfc ;
            rom[16564] = 8'h03 ;
            rom[16565] = 8'hf5 ;
            rom[16566] = 8'hca ;
            rom[16567] = 8'hd0 ;
            rom[16568] = 8'hee ;
            rom[16569] = 8'h0e ;
            rom[16570] = 8'h1b ;
            rom[16571] = 8'h0a ;
            rom[16572] = 8'hb8 ;
            rom[16573] = 8'he3 ;
            rom[16574] = 8'hca ;
            rom[16575] = 8'he3 ;
            rom[16576] = 8'h26 ;
            rom[16577] = 8'heb ;
            rom[16578] = 8'h1a ;
            rom[16579] = 8'hc5 ;
            rom[16580] = 8'h1d ;
            rom[16581] = 8'hf8 ;
            rom[16582] = 8'hd1 ;
            rom[16583] = 8'hd2 ;
            rom[16584] = 8'h05 ;
            rom[16585] = 8'hf0 ;
            rom[16586] = 8'hfc ;
            rom[16587] = 8'h09 ;
            rom[16588] = 8'he3 ;
            rom[16589] = 8'he9 ;
            rom[16590] = 8'h0f ;
            rom[16591] = 8'hff ;
            rom[16592] = 8'he4 ;
            rom[16593] = 8'hed ;
            rom[16594] = 8'hd1 ;
            rom[16595] = 8'hf1 ;
            rom[16596] = 8'hdb ;
            rom[16597] = 8'he7 ;
            rom[16598] = 8'h00 ;
            rom[16599] = 8'he2 ;
            rom[16600] = 8'h18 ;
            rom[16601] = 8'hf2 ;
            rom[16602] = 8'h27 ;
            rom[16603] = 8'h04 ;
            rom[16604] = 8'hc0 ;
            rom[16605] = 8'hf3 ;
            rom[16606] = 8'h13 ;
            rom[16607] = 8'hd7 ;
            rom[16608] = 8'h20 ;
            rom[16609] = 8'he0 ;
            rom[16610] = 8'h22 ;
            rom[16611] = 8'hf0 ;
            rom[16612] = 8'hfd ;
            rom[16613] = 8'hd0 ;
            rom[16614] = 8'hc4 ;
            rom[16615] = 8'hf5 ;
            rom[16616] = 8'hef ;
            rom[16617] = 8'he3 ;
            rom[16618] = 8'he0 ;
            rom[16619] = 8'h07 ;
            rom[16620] = 8'hf7 ;
            rom[16621] = 8'h1d ;
            rom[16622] = 8'h26 ;
            rom[16623] = 8'h13 ;
            rom[16624] = 8'hea ;
            rom[16625] = 8'h14 ;
            rom[16626] = 8'hfd ;
            rom[16627] = 8'hd7 ;
            rom[16628] = 8'he1 ;
            rom[16629] = 8'h0a ;
            rom[16630] = 8'h18 ;
            rom[16631] = 8'h17 ;
            rom[16632] = 8'h08 ;
            rom[16633] = 8'h1d ;
            rom[16634] = 8'h08 ;
            rom[16635] = 8'he4 ;
            rom[16636] = 8'hde ;
            rom[16637] = 8'hc6 ;
            rom[16638] = 8'hff ;
            rom[16639] = 8'hd8 ;
            rom[16640] = 8'hff ;
            rom[16641] = 8'hfa ;
            rom[16642] = 8'hfc ;
            rom[16643] = 8'h1b ;
            rom[16644] = 8'hec ;
            rom[16645] = 8'hdf ;
            rom[16646] = 8'h26 ;
            rom[16647] = 8'he7 ;
            rom[16648] = 8'hfe ;
            rom[16649] = 8'hfd ;
            rom[16650] = 8'h07 ;
            rom[16651] = 8'hdf ;
            rom[16652] = 8'hf7 ;
            rom[16653] = 8'h04 ;
            rom[16654] = 8'h0a ;
            rom[16655] = 8'hec ;
            rom[16656] = 8'h00 ;
            rom[16657] = 8'h08 ;
            rom[16658] = 8'h01 ;
            rom[16659] = 8'hef ;
            rom[16660] = 8'h34 ;
            rom[16661] = 8'he3 ;
            rom[16662] = 8'hca ;
            rom[16663] = 8'he8 ;
            rom[16664] = 8'h14 ;
            rom[16665] = 8'h18 ;
            rom[16666] = 8'h0a ;
            rom[16667] = 8'hfb ;
            rom[16668] = 8'he9 ;
            rom[16669] = 8'hff ;
            rom[16670] = 8'hfd ;
            rom[16671] = 8'hf1 ;
            rom[16672] = 8'h22 ;
            rom[16673] = 8'hc2 ;
            rom[16674] = 8'h16 ;
            rom[16675] = 8'h0d ;
            rom[16676] = 8'hec ;
            rom[16677] = 8'h22 ;
            rom[16678] = 8'hf9 ;
            rom[16679] = 8'h00 ;
            rom[16680] = 8'hd2 ;
            rom[16681] = 8'h10 ;
            rom[16682] = 8'heb ;
            rom[16683] = 8'hf1 ;
            rom[16684] = 8'h0f ;
            rom[16685] = 8'h43 ;
            rom[16686] = 8'hf4 ;
            rom[16687] = 8'h12 ;
            rom[16688] = 8'h0a ;
            rom[16689] = 8'h1e ;
            rom[16690] = 8'he3 ;
            rom[16691] = 8'hb8 ;
            rom[16692] = 8'h0a ;
            rom[16693] = 8'he6 ;
            rom[16694] = 8'hbb ;
            rom[16695] = 8'h1f ;
            rom[16696] = 8'h24 ;
            rom[16697] = 8'h0c ;
            rom[16698] = 8'hff ;
            rom[16699] = 8'he5 ;
            rom[16700] = 8'h1a ;
            rom[16701] = 8'he6 ;
            rom[16702] = 8'he3 ;
            rom[16703] = 8'he3 ;
            rom[16704] = 8'hf3 ;
            rom[16705] = 8'h14 ;
            rom[16706] = 8'hfd ;
            rom[16707] = 8'h14 ;
            rom[16708] = 8'h14 ;
            rom[16709] = 8'h10 ;
            rom[16710] = 8'hf7 ;
            rom[16711] = 8'h03 ;
            rom[16712] = 8'h11 ;
            rom[16713] = 8'h07 ;
            rom[16714] = 8'hf0 ;
            rom[16715] = 8'h06 ;
            rom[16716] = 8'h08 ;
            rom[16717] = 8'hfb ;
            rom[16718] = 8'hfc ;
            rom[16719] = 8'h28 ;
            rom[16720] = 8'he3 ;
            rom[16721] = 8'hb3 ;
            rom[16722] = 8'hf6 ;
            rom[16723] = 8'h12 ;
            rom[16724] = 8'hec ;
            rom[16725] = 8'h05 ;
            rom[16726] = 8'hde ;
            rom[16727] = 8'h0f ;
            rom[16728] = 8'h24 ;
            rom[16729] = 8'hea ;
            rom[16730] = 8'h25 ;
            rom[16731] = 8'h06 ;
            rom[16732] = 8'hf1 ;
            rom[16733] = 8'h0d ;
            rom[16734] = 8'h03 ;
            rom[16735] = 8'h13 ;
            rom[16736] = 8'h02 ;
            rom[16737] = 8'hde ;
            rom[16738] = 8'h03 ;
            rom[16739] = 8'hf3 ;
            rom[16740] = 8'hf0 ;
            rom[16741] = 8'h13 ;
            rom[16742] = 8'h00 ;
            rom[16743] = 8'hee ;
            rom[16744] = 8'hcd ;
            rom[16745] = 8'hd8 ;
            rom[16746] = 8'h1d ;
            rom[16747] = 8'hef ;
            rom[16748] = 8'h10 ;
            rom[16749] = 8'h06 ;
            rom[16750] = 8'h09 ;
            rom[16751] = 8'hed ;
            rom[16752] = 8'hf1 ;
            rom[16753] = 8'hcd ;
            rom[16754] = 8'h1e ;
            rom[16755] = 8'hde ;
            rom[16756] = 8'h03 ;
            rom[16757] = 8'h0e ;
            rom[16758] = 8'hf9 ;
            rom[16759] = 8'h21 ;
            rom[16760] = 8'hfb ;
            rom[16761] = 8'he7 ;
            rom[16762] = 8'hef ;
            rom[16763] = 8'hef ;
            rom[16764] = 8'hfc ;
            rom[16765] = 8'hf5 ;
            rom[16766] = 8'hd6 ;
            rom[16767] = 8'h00 ;
            rom[16768] = 8'hd6 ;
            rom[16769] = 8'h0a ;
            rom[16770] = 8'hfc ;
            rom[16771] = 8'h02 ;
            rom[16772] = 8'h0f ;
            rom[16773] = 8'hec ;
            rom[16774] = 8'h0f ;
            rom[16775] = 8'hf6 ;
            rom[16776] = 8'he2 ;
            rom[16777] = 8'hdc ;
            rom[16778] = 8'h39 ;
            rom[16779] = 8'h16 ;
            rom[16780] = 8'he5 ;
            rom[16781] = 8'hff ;
            rom[16782] = 8'hd7 ;
            rom[16783] = 8'h18 ;
            rom[16784] = 8'hff ;
            rom[16785] = 8'he1 ;
            rom[16786] = 8'hee ;
            rom[16787] = 8'he5 ;
            rom[16788] = 8'h23 ;
            rom[16789] = 8'hf2 ;
            rom[16790] = 8'hd5 ;
            rom[16791] = 8'h06 ;
            rom[16792] = 8'hfc ;
            rom[16793] = 8'h1a ;
            rom[16794] = 8'h1d ;
            rom[16795] = 8'hf9 ;
            rom[16796] = 8'h0f ;
            rom[16797] = 8'hf4 ;
            rom[16798] = 8'hec ;
            rom[16799] = 8'hec ;
            rom[16800] = 8'h1d ;
            rom[16801] = 8'h11 ;
            rom[16802] = 8'he0 ;
            rom[16803] = 8'h08 ;
            rom[16804] = 8'hf8 ;
            rom[16805] = 8'h08 ;
            rom[16806] = 8'he8 ;
            rom[16807] = 8'h16 ;
            rom[16808] = 8'h08 ;
            rom[16809] = 8'h00 ;
            rom[16810] = 8'h00 ;
            rom[16811] = 8'h02 ;
            rom[16812] = 8'h10 ;
            rom[16813] = 8'h1d ;
            rom[16814] = 8'hf3 ;
            rom[16815] = 8'he5 ;
            rom[16816] = 8'h13 ;
            rom[16817] = 8'hfe ;
            rom[16818] = 8'h02 ;
            rom[16819] = 8'he3 ;
            rom[16820] = 8'h09 ;
            rom[16821] = 8'hfa ;
            rom[16822] = 8'hfd ;
            rom[16823] = 8'hed ;
            rom[16824] = 8'hfe ;
            rom[16825] = 8'hff ;
            rom[16826] = 8'hff ;
            rom[16827] = 8'he0 ;
            rom[16828] = 8'h0b ;
            rom[16829] = 8'hf5 ;
            rom[16830] = 8'h0b ;
            rom[16831] = 8'hf2 ;
            rom[16832] = 8'hd3 ;
            rom[16833] = 8'he4 ;
            rom[16834] = 8'hea ;
            rom[16835] = 8'hfd ;
            rom[16836] = 8'hcf ;
            rom[16837] = 8'h13 ;
            rom[16838] = 8'hd9 ;
            rom[16839] = 8'h0c ;
            rom[16840] = 8'hbe ;
            rom[16841] = 8'hf2 ;
            rom[16842] = 8'h21 ;
            rom[16843] = 8'hfe ;
            rom[16844] = 8'hff ;
            rom[16845] = 8'hdd ;
            rom[16846] = 8'hf8 ;
            rom[16847] = 8'hf7 ;
            rom[16848] = 8'hfb ;
            rom[16849] = 8'he8 ;
            rom[16850] = 8'h04 ;
            rom[16851] = 8'hf1 ;
            rom[16852] = 8'he5 ;
            rom[16853] = 8'hf5 ;
            rom[16854] = 8'hf0 ;
            rom[16855] = 8'hf4 ;
            rom[16856] = 8'he9 ;
            rom[16857] = 8'hff ;
            rom[16858] = 8'h03 ;
            rom[16859] = 8'hf4 ;
            rom[16860] = 8'he8 ;
            rom[16861] = 8'he6 ;
            rom[16862] = 8'h01 ;
            rom[16863] = 8'h0c ;
            rom[16864] = 8'hc8 ;
            rom[16865] = 8'h10 ;
            rom[16866] = 8'hea ;
            rom[16867] = 8'hf5 ;
            rom[16868] = 8'h0b ;
            rom[16869] = 8'h19 ;
            rom[16870] = 8'h1d ;
            rom[16871] = 8'h10 ;
            rom[16872] = 8'h0b ;
            rom[16873] = 8'h0c ;
            rom[16874] = 8'hf9 ;
            rom[16875] = 8'he8 ;
            rom[16876] = 8'hfc ;
            rom[16877] = 8'he4 ;
            rom[16878] = 8'hdb ;
            rom[16879] = 8'h07 ;
            rom[16880] = 8'h27 ;
            rom[16881] = 8'hf8 ;
            rom[16882] = 8'h2b ;
            rom[16883] = 8'he9 ;
            rom[16884] = 8'h0e ;
            rom[16885] = 8'h33 ;
            rom[16886] = 8'hf4 ;
            rom[16887] = 8'hed ;
            rom[16888] = 8'hec ;
            rom[16889] = 8'he0 ;
            rom[16890] = 8'h14 ;
            rom[16891] = 8'hf2 ;
            rom[16892] = 8'h03 ;
            rom[16893] = 8'h16 ;
            rom[16894] = 8'h0e ;
            rom[16895] = 8'h12 ;
            rom[16896] = 8'hf4 ;
            rom[16897] = 8'h0d ;
            rom[16898] = 8'he6 ;
            rom[16899] = 8'hf1 ;
            rom[16900] = 8'h20 ;
            rom[16901] = 8'hfe ;
            rom[16902] = 8'hf3 ;
            rom[16903] = 8'hf5 ;
            rom[16904] = 8'hf9 ;
            rom[16905] = 8'h0b ;
            rom[16906] = 8'heb ;
            rom[16907] = 8'hf3 ;
            rom[16908] = 8'h11 ;
            rom[16909] = 8'h0f ;
            rom[16910] = 8'hff ;
            rom[16911] = 8'hf6 ;
            rom[16912] = 8'h01 ;
            rom[16913] = 8'h11 ;
            rom[16914] = 8'h0f ;
            rom[16915] = 8'hd3 ;
            rom[16916] = 8'h2e ;
            rom[16917] = 8'hf9 ;
            rom[16918] = 8'h1c ;
            rom[16919] = 8'h32 ;
            rom[16920] = 8'h06 ;
            rom[16921] = 8'h15 ;
            rom[16922] = 8'hdc ;
            rom[16923] = 8'hf8 ;
            rom[16924] = 8'hcb ;
            rom[16925] = 8'h15 ;
            rom[16926] = 8'h01 ;
            rom[16927] = 8'h0b ;
            rom[16928] = 8'h22 ;
            rom[16929] = 8'he6 ;
            rom[16930] = 8'hf1 ;
            rom[16931] = 8'hd0 ;
            rom[16932] = 8'hd1 ;
            rom[16933] = 8'hdb ;
            rom[16934] = 8'h21 ;
            rom[16935] = 8'hea ;
            rom[16936] = 8'hed ;
            rom[16937] = 8'hfc ;
            rom[16938] = 8'hf6 ;
            rom[16939] = 8'h1e ;
            rom[16940] = 8'h0b ;
            rom[16941] = 8'hef ;
            rom[16942] = 8'hf5 ;
            rom[16943] = 8'h17 ;
            rom[16944] = 8'hd6 ;
            rom[16945] = 8'hf6 ;
            rom[16946] = 8'hed ;
            rom[16947] = 8'hfd ;
            rom[16948] = 8'h09 ;
            rom[16949] = 8'h0f ;
            rom[16950] = 8'h0d ;
            rom[16951] = 8'he2 ;
            rom[16952] = 8'hec ;
            rom[16953] = 8'hfc ;
            rom[16954] = 8'h04 ;
            rom[16955] = 8'hdd ;
            rom[16956] = 8'hfa ;
            rom[16957] = 8'h02 ;
            rom[16958] = 8'h0e ;
            rom[16959] = 8'h1c ;
            rom[16960] = 8'h1f ;
            rom[16961] = 8'h1f ;
            rom[16962] = 8'h0c ;
            rom[16963] = 8'h07 ;
            rom[16964] = 8'h2c ;
            rom[16965] = 8'he4 ;
            rom[16966] = 8'he6 ;
            rom[16967] = 8'h0c ;
            rom[16968] = 8'h15 ;
            rom[16969] = 8'hdf ;
            rom[16970] = 8'hd7 ;
            rom[16971] = 8'he5 ;
            rom[16972] = 8'hf3 ;
            rom[16973] = 8'he6 ;
            rom[16974] = 8'hc9 ;
            rom[16975] = 8'h25 ;
            rom[16976] = 8'hc0 ;
            rom[16977] = 8'h13 ;
            rom[16978] = 8'hf4 ;
            rom[16979] = 8'hf9 ;
            rom[16980] = 8'hee ;
            rom[16981] = 8'h0f ;
            rom[16982] = 8'hf7 ;
            rom[16983] = 8'h24 ;
            rom[16984] = 8'hff ;
            rom[16985] = 8'he1 ;
            rom[16986] = 8'hff ;
            rom[16987] = 8'he8 ;
            rom[16988] = 8'h05 ;
            rom[16989] = 8'h04 ;
            rom[16990] = 8'h01 ;
            rom[16991] = 8'hf8 ;
            rom[16992] = 8'h0d ;
            rom[16993] = 8'h03 ;
            rom[16994] = 8'he9 ;
            rom[16995] = 8'hd8 ;
            rom[16996] = 8'he6 ;
            rom[16997] = 8'h03 ;
            rom[16998] = 8'hde ;
            rom[16999] = 8'h0d ;
            rom[17000] = 8'he7 ;
            rom[17001] = 8'hce ;
            rom[17002] = 8'h08 ;
            rom[17003] = 8'h29 ;
            rom[17004] = 8'hec ;
            rom[17005] = 8'he4 ;
            rom[17006] = 8'h1e ;
            rom[17007] = 8'h0f ;
            rom[17008] = 8'h0e ;
            rom[17009] = 8'hfb ;
            rom[17010] = 8'h14 ;
            rom[17011] = 8'h20 ;
            rom[17012] = 8'hdf ;
            rom[17013] = 8'he5 ;
            rom[17014] = 8'he2 ;
            rom[17015] = 8'h0a ;
            rom[17016] = 8'he7 ;
            rom[17017] = 8'h1a ;
            rom[17018] = 8'hae ;
            rom[17019] = 8'hf9 ;
            rom[17020] = 8'h10 ;
            rom[17021] = 8'h03 ;
            rom[17022] = 8'h08 ;
            rom[17023] = 8'h03 ;
            rom[17024] = 8'h28 ;
            rom[17025] = 8'hdc ;
            rom[17026] = 8'hd9 ;
            rom[17027] = 8'h05 ;
            rom[17028] = 8'hf5 ;
            rom[17029] = 8'hf3 ;
            rom[17030] = 8'hdf ;
            rom[17031] = 8'hf4 ;
            rom[17032] = 8'h1d ;
            rom[17033] = 8'hfd ;
            rom[17034] = 8'h09 ;
            rom[17035] = 8'hcb ;
            rom[17036] = 8'hf1 ;
            rom[17037] = 8'hf9 ;
            rom[17038] = 8'h08 ;
            rom[17039] = 8'h01 ;
            rom[17040] = 8'h09 ;
            rom[17041] = 8'hfe ;
            rom[17042] = 8'hd5 ;
            rom[17043] = 8'he1 ;
            rom[17044] = 8'he4 ;
            rom[17045] = 8'hf7 ;
            rom[17046] = 8'hdf ;
            rom[17047] = 8'hd3 ;
            rom[17048] = 8'hfd ;
            rom[17049] = 8'hfb ;
            rom[17050] = 8'h18 ;
            rom[17051] = 8'h01 ;
            rom[17052] = 8'h17 ;
            rom[17053] = 8'hc7 ;
            rom[17054] = 8'hed ;
            rom[17055] = 8'h04 ;
            rom[17056] = 8'hf4 ;
            rom[17057] = 8'h05 ;
            rom[17058] = 8'hbf ;
            rom[17059] = 8'hfc ;
            rom[17060] = 8'hf0 ;
            rom[17061] = 8'he7 ;
            rom[17062] = 8'he5 ;
            rom[17063] = 8'h11 ;
            rom[17064] = 8'h29 ;
            rom[17065] = 8'hf8 ;
            rom[17066] = 8'hec ;
            rom[17067] = 8'h12 ;
            rom[17068] = 8'h12 ;
            rom[17069] = 8'h08 ;
            rom[17070] = 8'he4 ;
            rom[17071] = 8'he0 ;
            rom[17072] = 8'h02 ;
            rom[17073] = 8'hea ;
            rom[17074] = 8'hfa ;
            rom[17075] = 8'hd1 ;
            rom[17076] = 8'h14 ;
            rom[17077] = 8'h00 ;
            rom[17078] = 8'hd4 ;
            rom[17079] = 8'hf4 ;
            rom[17080] = 8'h0c ;
            rom[17081] = 8'h09 ;
            rom[17082] = 8'h0c ;
            rom[17083] = 8'hf7 ;
            rom[17084] = 8'h0b ;
            rom[17085] = 8'he3 ;
            rom[17086] = 8'h11 ;
            rom[17087] = 8'he0 ;
            rom[17088] = 8'hf1 ;
            rom[17089] = 8'hdf ;
            rom[17090] = 8'hf6 ;
            rom[17091] = 8'h05 ;
            rom[17092] = 8'h17 ;
            rom[17093] = 8'hec ;
            rom[17094] = 8'he2 ;
            rom[17095] = 8'h01 ;
            rom[17096] = 8'h17 ;
            rom[17097] = 8'h1e ;
            rom[17098] = 8'h20 ;
            rom[17099] = 8'h37 ;
            rom[17100] = 8'h18 ;
            rom[17101] = 8'hef ;
            rom[17102] = 8'hf0 ;
            rom[17103] = 8'he1 ;
            rom[17104] = 8'hc8 ;
            rom[17105] = 8'h01 ;
            rom[17106] = 8'he6 ;
            rom[17107] = 8'heb ;
            rom[17108] = 8'hf8 ;
            rom[17109] = 8'he7 ;
            rom[17110] = 8'heb ;
            rom[17111] = 8'hf5 ;
            rom[17112] = 8'h10 ;
            rom[17113] = 8'hda ;
            rom[17114] = 8'h22 ;
            rom[17115] = 8'h13 ;
            rom[17116] = 8'hed ;
            rom[17117] = 8'h06 ;
            rom[17118] = 8'hf3 ;
            rom[17119] = 8'hf0 ;
            rom[17120] = 8'hf1 ;
            rom[17121] = 8'hfc ;
            rom[17122] = 8'h0e ;
            rom[17123] = 8'he8 ;
            rom[17124] = 8'h15 ;
            rom[17125] = 8'he9 ;
            rom[17126] = 8'h1f ;
            rom[17127] = 8'hbe ;
            rom[17128] = 8'hde ;
            rom[17129] = 8'h1a ;
            rom[17130] = 8'he7 ;
            rom[17131] = 8'hff ;
            rom[17132] = 8'hea ;
            rom[17133] = 8'h17 ;
            rom[17134] = 8'hee ;
            rom[17135] = 8'hf1 ;
            rom[17136] = 8'hee ;
            rom[17137] = 8'h2e ;
            rom[17138] = 8'hfa ;
            rom[17139] = 8'h07 ;
            rom[17140] = 8'hf4 ;
            rom[17141] = 8'he5 ;
            rom[17142] = 8'h20 ;
            rom[17143] = 8'h10 ;
            rom[17144] = 8'hd2 ;
            rom[17145] = 8'h14 ;
            rom[17146] = 8'h1f ;
            rom[17147] = 8'hfc ;
            rom[17148] = 8'hec ;
            rom[17149] = 8'hdd ;
            rom[17150] = 8'he9 ;
            rom[17151] = 8'he0 ;
            rom[17152] = 8'h0c ;
            rom[17153] = 8'hec ;
            rom[17154] = 8'h12 ;
            rom[17155] = 8'h1a ;
            rom[17156] = 8'hf0 ;
            rom[17157] = 8'h21 ;
            rom[17158] = 8'hbf ;
            rom[17159] = 8'hf7 ;
            rom[17160] = 8'hf6 ;
            rom[17161] = 8'h16 ;
            rom[17162] = 8'h0f ;
            rom[17163] = 8'h02 ;
            rom[17164] = 8'hf3 ;
            rom[17165] = 8'h14 ;
            rom[17166] = 8'h1f ;
            rom[17167] = 8'he8 ;
            rom[17168] = 8'h20 ;
            rom[17169] = 8'hf8 ;
            rom[17170] = 8'h08 ;
            rom[17171] = 8'h14 ;
            rom[17172] = 8'h14 ;
            rom[17173] = 8'hd9 ;
            rom[17174] = 8'h18 ;
            rom[17175] = 8'h01 ;
            rom[17176] = 8'hdb ;
            rom[17177] = 8'h1a ;
            rom[17178] = 8'h11 ;
            rom[17179] = 8'hc3 ;
            rom[17180] = 8'hfe ;
            rom[17181] = 8'h0a ;
            rom[17182] = 8'he3 ;
            rom[17183] = 8'h09 ;
            rom[17184] = 8'hd5 ;
            rom[17185] = 8'he0 ;
            rom[17186] = 8'h11 ;
            rom[17187] = 8'hc3 ;
            rom[17188] = 8'hf8 ;
            rom[17189] = 8'hf5 ;
            rom[17190] = 8'h03 ;
            rom[17191] = 8'hc5 ;
            rom[17192] = 8'h0a ;
            rom[17193] = 8'hc4 ;
            rom[17194] = 8'h07 ;
            rom[17195] = 8'hfb ;
            rom[17196] = 8'h12 ;
            rom[17197] = 8'h11 ;
            rom[17198] = 8'he1 ;
            rom[17199] = 8'hf9 ;
            rom[17200] = 8'hf7 ;
            rom[17201] = 8'hf1 ;
            rom[17202] = 8'h05 ;
            rom[17203] = 8'hd6 ;
            rom[17204] = 8'h1e ;
            rom[17205] = 8'he2 ;
            rom[17206] = 8'h0f ;
            rom[17207] = 8'he7 ;
            rom[17208] = 8'h02 ;
            rom[17209] = 8'hde ;
            rom[17210] = 8'hea ;
            rom[17211] = 8'h0a ;
            rom[17212] = 8'hed ;
            rom[17213] = 8'hf6 ;
            rom[17214] = 8'h05 ;
            rom[17215] = 8'h06 ;
            rom[17216] = 8'he7 ;
            rom[17217] = 8'hfb ;
            rom[17218] = 8'h02 ;
            rom[17219] = 8'hd5 ;
            rom[17220] = 8'h00 ;
            rom[17221] = 8'hd6 ;
            rom[17222] = 8'hef ;
            rom[17223] = 8'h02 ;
            rom[17224] = 8'h0a ;
            rom[17225] = 8'hfe ;
            rom[17226] = 8'he9 ;
            rom[17227] = 8'h23 ;
            rom[17228] = 8'hd9 ;
            rom[17229] = 8'h06 ;
            rom[17230] = 8'h03 ;
            rom[17231] = 8'h00 ;
            rom[17232] = 8'hd4 ;
            rom[17233] = 8'h0b ;
            rom[17234] = 8'hea ;
            rom[17235] = 8'h09 ;
            rom[17236] = 8'h0f ;
            rom[17237] = 8'h1e ;
            rom[17238] = 8'h07 ;
            rom[17239] = 8'hef ;
            rom[17240] = 8'h04 ;
            rom[17241] = 8'hd4 ;
            rom[17242] = 8'h20 ;
            rom[17243] = 8'h25 ;
            rom[17244] = 8'hd5 ;
            rom[17245] = 8'he0 ;
            rom[17246] = 8'h12 ;
            rom[17247] = 8'hf8 ;
            rom[17248] = 8'he1 ;
            rom[17249] = 8'h0a ;
            rom[17250] = 8'hd1 ;
            rom[17251] = 8'h09 ;
            rom[17252] = 8'hdf ;
            rom[17253] = 8'h03 ;
            rom[17254] = 8'hff ;
            rom[17255] = 8'hf7 ;
            rom[17256] = 8'hf0 ;
            rom[17257] = 8'hf3 ;
            rom[17258] = 8'h09 ;
            rom[17259] = 8'h00 ;
            rom[17260] = 8'h1d ;
            rom[17261] = 8'hf9 ;
            rom[17262] = 8'h06 ;
            rom[17263] = 8'hea ;
            rom[17264] = 8'hd1 ;
            rom[17265] = 8'he5 ;
            rom[17266] = 8'h23 ;
            rom[17267] = 8'h05 ;
            rom[17268] = 8'hcc ;
            rom[17269] = 8'hef ;
            rom[17270] = 8'he8 ;
            rom[17271] = 8'hfa ;
            rom[17272] = 8'hff ;
            rom[17273] = 8'hf5 ;
            rom[17274] = 8'hca ;
            rom[17275] = 8'he5 ;
            rom[17276] = 8'hde ;
            rom[17277] = 8'h00 ;
            rom[17278] = 8'hdb ;
            rom[17279] = 8'h0f ;
            rom[17280] = 8'h05 ;
            rom[17281] = 8'h14 ;
            rom[17282] = 8'hf9 ;
            rom[17283] = 8'h24 ;
            rom[17284] = 8'he6 ;
            rom[17285] = 8'h08 ;
            rom[17286] = 8'hf6 ;
            rom[17287] = 8'hda ;
            rom[17288] = 8'hfa ;
            rom[17289] = 8'hec ;
            rom[17290] = 8'h0d ;
            rom[17291] = 8'hf5 ;
            rom[17292] = 8'he7 ;
            rom[17293] = 8'hf1 ;
            rom[17294] = 8'hf2 ;
            rom[17295] = 8'h12 ;
            rom[17296] = 8'h0f ;
            rom[17297] = 8'h0d ;
            rom[17298] = 8'hf1 ;
            rom[17299] = 8'h01 ;
            rom[17300] = 8'hf9 ;
            rom[17301] = 8'h08 ;
            rom[17302] = 8'h11 ;
            rom[17303] = 8'he2 ;
            rom[17304] = 8'h23 ;
            rom[17305] = 8'hee ;
            rom[17306] = 8'h03 ;
            rom[17307] = 8'hef ;
            rom[17308] = 8'hd7 ;
            rom[17309] = 8'hf9 ;
            rom[17310] = 8'h12 ;
            rom[17311] = 8'h0e ;
            rom[17312] = 8'he1 ;
            rom[17313] = 8'h12 ;
            rom[17314] = 8'hf5 ;
            rom[17315] = 8'hf8 ;
            rom[17316] = 8'h06 ;
            rom[17317] = 8'he0 ;
            rom[17318] = 8'hfc ;
            rom[17319] = 8'hea ;
            rom[17320] = 8'h01 ;
            rom[17321] = 8'hd6 ;
            rom[17322] = 8'hfd ;
            rom[17323] = 8'h25 ;
            rom[17324] = 8'h03 ;
            rom[17325] = 8'hf1 ;
            rom[17326] = 8'he4 ;
            rom[17327] = 8'hff ;
            rom[17328] = 8'h0a ;
            rom[17329] = 8'h0b ;
            rom[17330] = 8'heb ;
            rom[17331] = 8'h16 ;
            rom[17332] = 8'hdc ;
            rom[17333] = 8'h01 ;
            rom[17334] = 8'h1b ;
            rom[17335] = 8'hf5 ;
            rom[17336] = 8'h21 ;
            rom[17337] = 8'hf8 ;
            rom[17338] = 8'hef ;
            rom[17339] = 8'hec ;
            rom[17340] = 8'hfe ;
            rom[17341] = 8'h06 ;
            rom[17342] = 8'hfb ;
            rom[17343] = 8'h05 ;
            rom[17344] = 8'h1e ;
            rom[17345] = 8'h0a ;
            rom[17346] = 8'h0c ;
            rom[17347] = 8'hdd ;
            rom[17348] = 8'he3 ;
            rom[17349] = 8'hde ;
            rom[17350] = 8'hce ;
            rom[17351] = 8'h00 ;
            rom[17352] = 8'h01 ;
            rom[17353] = 8'hed ;
            rom[17354] = 8'hde ;
            rom[17355] = 8'hc6 ;
            rom[17356] = 8'h00 ;
            rom[17357] = 8'hf7 ;
            rom[17358] = 8'he7 ;
            rom[17359] = 8'h10 ;
            rom[17360] = 8'h0d ;
            rom[17361] = 8'h04 ;
            rom[17362] = 8'h07 ;
            rom[17363] = 8'hf2 ;
            rom[17364] = 8'heb ;
            rom[17365] = 8'he7 ;
            rom[17366] = 8'he3 ;
            rom[17367] = 8'h1b ;
            rom[17368] = 8'h11 ;
            rom[17369] = 8'h03 ;
            rom[17370] = 8'hfa ;
            rom[17371] = 8'h0d ;
            rom[17372] = 8'hd5 ;
            rom[17373] = 8'h2f ;
            rom[17374] = 8'hee ;
            rom[17375] = 8'hcf ;
            rom[17376] = 8'h30 ;
            rom[17377] = 8'h14 ;
            rom[17378] = 8'hff ;
            rom[17379] = 8'h0e ;
            rom[17380] = 8'hdc ;
            rom[17381] = 8'h10 ;
            rom[17382] = 8'hde ;
            rom[17383] = 8'hdb ;
            rom[17384] = 8'h12 ;
            rom[17385] = 8'h05 ;
            rom[17386] = 8'heb ;
            rom[17387] = 8'hff ;
            rom[17388] = 8'hf3 ;
            rom[17389] = 8'he9 ;
            rom[17390] = 8'h24 ;
            rom[17391] = 8'h22 ;
            rom[17392] = 8'h0f ;
            rom[17393] = 8'he0 ;
            rom[17394] = 8'hd5 ;
            rom[17395] = 8'h0f ;
            rom[17396] = 8'he3 ;
            rom[17397] = 8'he7 ;
            rom[17398] = 8'hd4 ;
            rom[17399] = 8'h0d ;
            rom[17400] = 8'hf2 ;
            rom[17401] = 8'hf1 ;
            rom[17402] = 8'he3 ;
            rom[17403] = 8'hf5 ;
            rom[17404] = 8'hf0 ;
            rom[17405] = 8'h01 ;
            rom[17406] = 8'hfe ;
            rom[17407] = 8'h0d ;
            rom[17408] = 8'hed ;
            rom[17409] = 8'h04 ;
            rom[17410] = 8'he8 ;
            rom[17411] = 8'hea ;
            rom[17412] = 8'hf5 ;
            rom[17413] = 8'hfb ;
            rom[17414] = 8'hed ;
            rom[17415] = 8'hdc ;
            rom[17416] = 8'h0b ;
            rom[17417] = 8'h1e ;
            rom[17418] = 8'h1e ;
            rom[17419] = 8'h13 ;
            rom[17420] = 8'h0d ;
            rom[17421] = 8'h17 ;
            rom[17422] = 8'h00 ;
            rom[17423] = 8'hbf ;
            rom[17424] = 8'hfe ;
            rom[17425] = 8'heb ;
            rom[17426] = 8'h1c ;
            rom[17427] = 8'hea ;
            rom[17428] = 8'hff ;
            rom[17429] = 8'hdb ;
            rom[17430] = 8'h02 ;
            rom[17431] = 8'hf6 ;
            rom[17432] = 8'hd9 ;
            rom[17433] = 8'h0f ;
            rom[17434] = 8'hd2 ;
            rom[17435] = 8'hcc ;
            rom[17436] = 8'he0 ;
            rom[17437] = 8'hde ;
            rom[17438] = 8'hf5 ;
            rom[17439] = 8'hfb ;
            rom[17440] = 8'hd7 ;
            rom[17441] = 8'hea ;
            rom[17442] = 8'hd7 ;
            rom[17443] = 8'hf3 ;
            rom[17444] = 8'h21 ;
            rom[17445] = 8'hc8 ;
            rom[17446] = 8'hf9 ;
            rom[17447] = 8'hec ;
            rom[17448] = 8'hef ;
            rom[17449] = 8'h06 ;
            rom[17450] = 8'hf5 ;
            rom[17451] = 8'hfc ;
            rom[17452] = 8'hfd ;
            rom[17453] = 8'h09 ;
            rom[17454] = 8'h04 ;
            rom[17455] = 8'hfe ;
            rom[17456] = 8'he9 ;
            rom[17457] = 8'hf5 ;
            rom[17458] = 8'hf3 ;
            rom[17459] = 8'hf7 ;
            rom[17460] = 8'hf7 ;
            rom[17461] = 8'h00 ;
            rom[17462] = 8'hd8 ;
            rom[17463] = 8'he4 ;
            rom[17464] = 8'hc9 ;
            rom[17465] = 8'h08 ;
            rom[17466] = 8'he2 ;
            rom[17467] = 8'hf5 ;
            rom[17468] = 8'hc5 ;
            rom[17469] = 8'hff ;
            rom[17470] = 8'hf4 ;
            rom[17471] = 8'hf6 ;
            rom[17472] = 8'h12 ;
            rom[17473] = 8'hf3 ;
            rom[17474] = 8'h10 ;
            rom[17475] = 8'hf3 ;
            rom[17476] = 8'h0f ;
            rom[17477] = 8'hf0 ;
            rom[17478] = 8'hdd ;
            rom[17479] = 8'hf2 ;
            rom[17480] = 8'h18 ;
            rom[17481] = 8'h08 ;
            rom[17482] = 8'h0c ;
            rom[17483] = 8'h05 ;
            rom[17484] = 8'hc1 ;
            rom[17485] = 8'h00 ;
            rom[17486] = 8'h0a ;
            rom[17487] = 8'hf3 ;
            rom[17488] = 8'hee ;
            rom[17489] = 8'hfe ;
            rom[17490] = 8'h0b ;
            rom[17491] = 8'hf5 ;
            rom[17492] = 8'he5 ;
            rom[17493] = 8'h00 ;
            rom[17494] = 8'h10 ;
            rom[17495] = 8'h17 ;
            rom[17496] = 8'hfa ;
            rom[17497] = 8'hd4 ;
            rom[17498] = 8'h06 ;
            rom[17499] = 8'h03 ;
            rom[17500] = 8'hdb ;
            rom[17501] = 8'hec ;
            rom[17502] = 8'h0e ;
            rom[17503] = 8'hf8 ;
            rom[17504] = 8'hf2 ;
            rom[17505] = 8'hf8 ;
            rom[17506] = 8'hf2 ;
            rom[17507] = 8'hcf ;
            rom[17508] = 8'he2 ;
            rom[17509] = 8'h17 ;
            rom[17510] = 8'h02 ;
            rom[17511] = 8'hdb ;
            rom[17512] = 8'he1 ;
            rom[17513] = 8'hec ;
            rom[17514] = 8'hfc ;
            rom[17515] = 8'h02 ;
            rom[17516] = 8'h02 ;
            rom[17517] = 8'hc2 ;
            rom[17518] = 8'h12 ;
            rom[17519] = 8'h03 ;
            rom[17520] = 8'h01 ;
            rom[17521] = 8'he3 ;
            rom[17522] = 8'h20 ;
            rom[17523] = 8'hed ;
            rom[17524] = 8'hf5 ;
            rom[17525] = 8'hff ;
            rom[17526] = 8'he3 ;
            rom[17527] = 8'hfc ;
            rom[17528] = 8'h0e ;
            rom[17529] = 8'h17 ;
            rom[17530] = 8'he5 ;
            rom[17531] = 8'hf9 ;
            rom[17532] = 8'hff ;
            rom[17533] = 8'hf0 ;
            rom[17534] = 8'hce ;
            rom[17535] = 8'hf4 ;
            rom[17536] = 8'hd9 ;
            rom[17537] = 8'he4 ;
            rom[17538] = 8'h21 ;
            rom[17539] = 8'hf8 ;
            rom[17540] = 8'h07 ;
            rom[17541] = 8'hfd ;
            rom[17542] = 8'hf6 ;
            rom[17543] = 8'hd7 ;
            rom[17544] = 8'h07 ;
            rom[17545] = 8'h21 ;
            rom[17546] = 8'h1e ;
            rom[17547] = 8'h14 ;
            rom[17548] = 8'hbb ;
            rom[17549] = 8'h21 ;
            rom[17550] = 8'h22 ;
            rom[17551] = 8'h07 ;
            rom[17552] = 8'h2c ;
            rom[17553] = 8'he6 ;
            rom[17554] = 8'hdf ;
            rom[17555] = 8'hf0 ;
            rom[17556] = 8'h17 ;
            rom[17557] = 8'he4 ;
            rom[17558] = 8'hdf ;
            rom[17559] = 8'h0b ;
            rom[17560] = 8'hcf ;
            rom[17561] = 8'he8 ;
            rom[17562] = 8'hfb ;
            rom[17563] = 8'hcd ;
            rom[17564] = 8'he5 ;
            rom[17565] = 8'h29 ;
            rom[17566] = 8'he6 ;
            rom[17567] = 8'h02 ;
            rom[17568] = 8'h03 ;
            rom[17569] = 8'hf2 ;
            rom[17570] = 8'hfe ;
            rom[17571] = 8'hf9 ;
            rom[17572] = 8'h0f ;
            rom[17573] = 8'h10 ;
            rom[17574] = 8'h06 ;
            rom[17575] = 8'hde ;
            rom[17576] = 8'h00 ;
            rom[17577] = 8'hce ;
            rom[17578] = 8'h13 ;
            rom[17579] = 8'h1e ;
            rom[17580] = 8'h07 ;
            rom[17581] = 8'h03 ;
            rom[17582] = 8'h21 ;
            rom[17583] = 8'he1 ;
            rom[17584] = 8'hf9 ;
            rom[17585] = 8'hc1 ;
            rom[17586] = 8'he2 ;
            rom[17587] = 8'hf5 ;
            rom[17588] = 8'he9 ;
            rom[17589] = 8'hcc ;
            rom[17590] = 8'hfd ;
            rom[17591] = 8'hed ;
            rom[17592] = 8'h14 ;
            rom[17593] = 8'hd4 ;
            rom[17594] = 8'h1e ;
            rom[17595] = 8'h18 ;
            rom[17596] = 8'h01 ;
            rom[17597] = 8'hf6 ;
            rom[17598] = 8'h11 ;
            rom[17599] = 8'h08 ;
            rom[17600] = 8'hd7 ;
            rom[17601] = 8'hfd ;
            rom[17602] = 8'h1e ;
            rom[17603] = 8'he7 ;
            rom[17604] = 8'hfd ;
            rom[17605] = 8'hfa ;
            rom[17606] = 8'h2b ;
            rom[17607] = 8'h07 ;
            rom[17608] = 8'he6 ;
            rom[17609] = 8'h24 ;
            rom[17610] = 8'he4 ;
            rom[17611] = 8'h21 ;
            rom[17612] = 8'he5 ;
            rom[17613] = 8'hda ;
            rom[17614] = 8'h15 ;
            rom[17615] = 8'hea ;
            rom[17616] = 8'h12 ;
            rom[17617] = 8'h22 ;
            rom[17618] = 8'hf1 ;
            rom[17619] = 8'hc2 ;
            rom[17620] = 8'hf7 ;
            rom[17621] = 8'h2f ;
            rom[17622] = 8'h20 ;
            rom[17623] = 8'hed ;
            rom[17624] = 8'h43 ;
            rom[17625] = 8'he4 ;
            rom[17626] = 8'h07 ;
            rom[17627] = 8'hde ;
            rom[17628] = 8'hac ;
            rom[17629] = 8'hff ;
            rom[17630] = 8'hf7 ;
            rom[17631] = 8'h03 ;
            rom[17632] = 8'he9 ;
            rom[17633] = 8'h12 ;
            rom[17634] = 8'h0a ;
            rom[17635] = 8'hf2 ;
            rom[17636] = 8'he6 ;
            rom[17637] = 8'hdb ;
            rom[17638] = 8'he3 ;
            rom[17639] = 8'hf3 ;
            rom[17640] = 8'h1e ;
            rom[17641] = 8'hda ;
            rom[17642] = 8'h17 ;
            rom[17643] = 8'hff ;
            rom[17644] = 8'h21 ;
            rom[17645] = 8'hf8 ;
            rom[17646] = 8'hf1 ;
            rom[17647] = 8'hf5 ;
            rom[17648] = 8'he5 ;
            rom[17649] = 8'he2 ;
            rom[17650] = 8'hfc ;
            rom[17651] = 8'h0c ;
            rom[17652] = 8'hfa ;
            rom[17653] = 8'h19 ;
            rom[17654] = 8'h04 ;
            rom[17655] = 8'h07 ;
            rom[17656] = 8'hf8 ;
            rom[17657] = 8'h2f ;
            rom[17658] = 8'hd7 ;
            rom[17659] = 8'h04 ;
            rom[17660] = 8'h09 ;
            rom[17661] = 8'hf6 ;
            rom[17662] = 8'hdb ;
            rom[17663] = 8'hb9 ;
            rom[17664] = 8'hfa ;
            rom[17665] = 8'h22 ;
            rom[17666] = 8'hfa ;
            rom[17667] = 8'h04 ;
            rom[17668] = 8'h14 ;
            rom[17669] = 8'hff ;
            rom[17670] = 8'h06 ;
            rom[17671] = 8'hf1 ;
            rom[17672] = 8'h32 ;
            rom[17673] = 8'hee ;
            rom[17674] = 8'he7 ;
            rom[17675] = 8'hdb ;
            rom[17676] = 8'h04 ;
            rom[17677] = 8'hfe ;
            rom[17678] = 8'hf4 ;
            rom[17679] = 8'hf9 ;
            rom[17680] = 8'hfa ;
            rom[17681] = 8'h10 ;
            rom[17682] = 8'hf0 ;
            rom[17683] = 8'he5 ;
            rom[17684] = 8'hfd ;
            rom[17685] = 8'hfe ;
            rom[17686] = 8'h0b ;
            rom[17687] = 8'hfb ;
            rom[17688] = 8'h2a ;
            rom[17689] = 8'hed ;
            rom[17690] = 8'hee ;
            rom[17691] = 8'h08 ;
            rom[17692] = 8'hf2 ;
            rom[17693] = 8'h2f ;
            rom[17694] = 8'h14 ;
            rom[17695] = 8'hd2 ;
            rom[17696] = 8'hfb ;
            rom[17697] = 8'hcb ;
            rom[17698] = 8'h0e ;
            rom[17699] = 8'h00 ;
            rom[17700] = 8'he9 ;
            rom[17701] = 8'hee ;
            rom[17702] = 8'h27 ;
            rom[17703] = 8'h18 ;
            rom[17704] = 8'h08 ;
            rom[17705] = 8'he7 ;
            rom[17706] = 8'hfb ;
            rom[17707] = 8'h01 ;
            rom[17708] = 8'h17 ;
            rom[17709] = 8'hf2 ;
            rom[17710] = 8'h19 ;
            rom[17711] = 8'he7 ;
            rom[17712] = 8'he9 ;
            rom[17713] = 8'h1b ;
            rom[17714] = 8'h19 ;
            rom[17715] = 8'he9 ;
            rom[17716] = 8'hef ;
            rom[17717] = 8'he3 ;
            rom[17718] = 8'h0f ;
            rom[17719] = 8'hfe ;
            rom[17720] = 8'h35 ;
            rom[17721] = 8'h16 ;
            rom[17722] = 8'hf0 ;
            rom[17723] = 8'hdb ;
            rom[17724] = 8'he7 ;
            rom[17725] = 8'hc4 ;
            rom[17726] = 8'h1f ;
            rom[17727] = 8'h0f ;
            rom[17728] = 8'h06 ;
            rom[17729] = 8'h0c ;
            rom[17730] = 8'h19 ;
            rom[17731] = 8'h14 ;
            rom[17732] = 8'h0d ;
            rom[17733] = 8'h1a ;
            rom[17734] = 8'he8 ;
            rom[17735] = 8'hf9 ;
            rom[17736] = 8'hf9 ;
            rom[17737] = 8'h03 ;
            rom[17738] = 8'hcd ;
            rom[17739] = 8'hf2 ;
            rom[17740] = 8'hd4 ;
            rom[17741] = 8'hba ;
            rom[17742] = 8'hf6 ;
            rom[17743] = 8'hf4 ;
            rom[17744] = 8'h31 ;
            rom[17745] = 8'h25 ;
            rom[17746] = 8'hfe ;
            rom[17747] = 8'h15 ;
            rom[17748] = 8'h0d ;
            rom[17749] = 8'h19 ;
            rom[17750] = 8'he2 ;
            rom[17751] = 8'hf0 ;
            rom[17752] = 8'h27 ;
            rom[17753] = 8'h01 ;
            rom[17754] = 8'he0 ;
            rom[17755] = 8'h04 ;
            rom[17756] = 8'h2a ;
            rom[17757] = 8'h0a ;
            rom[17758] = 8'hc3 ;
            rom[17759] = 8'hea ;
            rom[17760] = 8'h21 ;
            rom[17761] = 8'h0a ;
            rom[17762] = 8'h04 ;
            rom[17763] = 8'he9 ;
            rom[17764] = 8'hff ;
            rom[17765] = 8'hf1 ;
            rom[17766] = 8'hf2 ;
            rom[17767] = 8'h11 ;
            rom[17768] = 8'h37 ;
            rom[17769] = 8'hff ;
            rom[17770] = 8'h0c ;
            rom[17771] = 8'h0a ;
            rom[17772] = 8'hff ;
            rom[17773] = 8'h0a ;
            rom[17774] = 8'he9 ;
            rom[17775] = 8'h0c ;
            rom[17776] = 8'h0a ;
            rom[17777] = 8'hd1 ;
            rom[17778] = 8'h07 ;
            rom[17779] = 8'h2d ;
            rom[17780] = 8'h20 ;
            rom[17781] = 8'hf1 ;
            rom[17782] = 8'hf1 ;
            rom[17783] = 8'he6 ;
            rom[17784] = 8'h10 ;
            rom[17785] = 8'hfc ;
            rom[17786] = 8'hd7 ;
            rom[17787] = 8'hef ;
            rom[17788] = 8'h05 ;
            rom[17789] = 8'h16 ;
            rom[17790] = 8'h1f ;
            rom[17791] = 8'h17 ;
            rom[17792] = 8'hd3 ;
            rom[17793] = 8'hfe ;
            rom[17794] = 8'h06 ;
            rom[17795] = 8'h0c ;
            rom[17796] = 8'hec ;
            rom[17797] = 8'h05 ;
            rom[17798] = 8'h0d ;
            rom[17799] = 8'hf6 ;
            rom[17800] = 8'h25 ;
            rom[17801] = 8'hbc ;
            rom[17802] = 8'hfe ;
            rom[17803] = 8'hbb ;
            rom[17804] = 8'hfb ;
            rom[17805] = 8'h1d ;
            rom[17806] = 8'h02 ;
            rom[17807] = 8'hfa ;
            rom[17808] = 8'hb5 ;
            rom[17809] = 8'h0c ;
            rom[17810] = 8'h11 ;
            rom[17811] = 8'hd9 ;
            rom[17812] = 8'hd4 ;
            rom[17813] = 8'hdb ;
            rom[17814] = 8'h13 ;
            rom[17815] = 8'h1a ;
            rom[17816] = 8'h10 ;
            rom[17817] = 8'hf3 ;
            rom[17818] = 8'hec ;
            rom[17819] = 8'h0d ;
            rom[17820] = 8'h16 ;
            rom[17821] = 8'hdc ;
            rom[17822] = 8'h24 ;
            rom[17823] = 8'he5 ;
            rom[17824] = 8'he8 ;
            rom[17825] = 8'h06 ;
            rom[17826] = 8'hf4 ;
            rom[17827] = 8'hfd ;
            rom[17828] = 8'hcf ;
            rom[17829] = 8'h01 ;
            rom[17830] = 8'h29 ;
            rom[17831] = 8'h1a ;
            rom[17832] = 8'hf8 ;
            rom[17833] = 8'hf5 ;
            rom[17834] = 8'h06 ;
            rom[17835] = 8'h1b ;
            rom[17836] = 8'h02 ;
            rom[17837] = 8'hd6 ;
            rom[17838] = 8'h20 ;
            rom[17839] = 8'hf3 ;
            rom[17840] = 8'h18 ;
            rom[17841] = 8'h00 ;
            rom[17842] = 8'hd4 ;
            rom[17843] = 8'h0a ;
            rom[17844] = 8'hde ;
            rom[17845] = 8'hd3 ;
            rom[17846] = 8'h13 ;
            rom[17847] = 8'h2e ;
            rom[17848] = 8'h37 ;
            rom[17849] = 8'hd3 ;
            rom[17850] = 8'hff ;
            rom[17851] = 8'h0d ;
            rom[17852] = 8'h0e ;
            rom[17853] = 8'he1 ;
            rom[17854] = 8'h0e ;
            rom[17855] = 8'h13 ;
            rom[17856] = 8'h08 ;
            rom[17857] = 8'hed ;
            rom[17858] = 8'hce ;
            rom[17859] = 8'hed ;
            rom[17860] = 8'hfa ;
            rom[17861] = 8'he9 ;
            rom[17862] = 8'he1 ;
            rom[17863] = 8'hb8 ;
            rom[17864] = 8'hf4 ;
            rom[17865] = 8'hd9 ;
            rom[17866] = 8'he6 ;
            rom[17867] = 8'he4 ;
            rom[17868] = 8'he4 ;
            rom[17869] = 8'h00 ;
            rom[17870] = 8'hcf ;
            rom[17871] = 8'h24 ;
            rom[17872] = 8'h15 ;
            rom[17873] = 8'h1d ;
            rom[17874] = 8'h0b ;
            rom[17875] = 8'h03 ;
            rom[17876] = 8'hff ;
            rom[17877] = 8'hfe ;
            rom[17878] = 8'hf0 ;
            rom[17879] = 8'h00 ;
            rom[17880] = 8'he6 ;
            rom[17881] = 8'hff ;
            rom[17882] = 8'hc8 ;
            rom[17883] = 8'h14 ;
            rom[17884] = 8'he6 ;
            rom[17885] = 8'h1b ;
            rom[17886] = 8'hc0 ;
            rom[17887] = 8'h05 ;
            rom[17888] = 8'h0d ;
            rom[17889] = 8'h00 ;
            rom[17890] = 8'he5 ;
            rom[17891] = 8'h10 ;
            rom[17892] = 8'h10 ;
            rom[17893] = 8'hec ;
            rom[17894] = 8'h05 ;
            rom[17895] = 8'h0d ;
            rom[17896] = 8'he9 ;
            rom[17897] = 8'hcf ;
            rom[17898] = 8'he7 ;
            rom[17899] = 8'hf8 ;
            rom[17900] = 8'hf3 ;
            rom[17901] = 8'he9 ;
            rom[17902] = 8'h0d ;
            rom[17903] = 8'h22 ;
            rom[17904] = 8'h0c ;
            rom[17905] = 8'h02 ;
            rom[17906] = 8'h07 ;
            rom[17907] = 8'h1b ;
            rom[17908] = 8'h2a ;
            rom[17909] = 8'h1a ;
            rom[17910] = 8'he4 ;
            rom[17911] = 8'hc8 ;
            rom[17912] = 8'he6 ;
            rom[17913] = 8'hf3 ;
            rom[17914] = 8'hd9 ;
            rom[17915] = 8'h25 ;
            rom[17916] = 8'h1b ;
            rom[17917] = 8'hfb ;
            rom[17918] = 8'h0a ;
            rom[17919] = 8'he8 ;
            rom[17920] = 8'hca ;
            rom[17921] = 8'h01 ;
            rom[17922] = 8'h03 ;
            rom[17923] = 8'hee ;
            rom[17924] = 8'hf9 ;
            rom[17925] = 8'h18 ;
            rom[17926] = 8'hf2 ;
            rom[17927] = 8'hf3 ;
            rom[17928] = 8'hff ;
            rom[17929] = 8'hf2 ;
            rom[17930] = 8'h04 ;
            rom[17931] = 8'h05 ;
            rom[17932] = 8'h35 ;
            rom[17933] = 8'h2b ;
            rom[17934] = 8'h27 ;
            rom[17935] = 8'hf5 ;
            rom[17936] = 8'hf9 ;
            rom[17937] = 8'heb ;
            rom[17938] = 8'hf5 ;
            rom[17939] = 8'hf4 ;
            rom[17940] = 8'hfb ;
            rom[17941] = 8'hf1 ;
            rom[17942] = 8'h07 ;
            rom[17943] = 8'h02 ;
            rom[17944] = 8'h18 ;
            rom[17945] = 8'h13 ;
            rom[17946] = 8'h13 ;
            rom[17947] = 8'h0f ;
            rom[17948] = 8'h0f ;
            rom[17949] = 8'hf1 ;
            rom[17950] = 8'h10 ;
            rom[17951] = 8'he8 ;
            rom[17952] = 8'hfc ;
            rom[17953] = 8'hfa ;
            rom[17954] = 8'h10 ;
            rom[17955] = 8'he6 ;
            rom[17956] = 8'hd8 ;
            rom[17957] = 8'h0e ;
            rom[17958] = 8'h0f ;
            rom[17959] = 8'h0c ;
            rom[17960] = 8'h21 ;
            rom[17961] = 8'h07 ;
            rom[17962] = 8'h16 ;
            rom[17963] = 8'h10 ;
            rom[17964] = 8'h11 ;
            rom[17965] = 8'h07 ;
            rom[17966] = 8'hd8 ;
            rom[17967] = 8'hc6 ;
            rom[17968] = 8'hf9 ;
            rom[17969] = 8'h17 ;
            rom[17970] = 8'h23 ;
            rom[17971] = 8'hdb ;
            rom[17972] = 8'he7 ;
            rom[17973] = 8'he4 ;
            rom[17974] = 8'h06 ;
            rom[17975] = 8'h1c ;
            rom[17976] = 8'h0c ;
            rom[17977] = 8'hf7 ;
            rom[17978] = 8'hfd ;
            rom[17979] = 8'hf9 ;
            rom[17980] = 8'hfb ;
            rom[17981] = 8'hfe ;
            rom[17982] = 8'h02 ;
            rom[17983] = 8'hf8 ;
            rom[17984] = 8'h16 ;
            rom[17985] = 8'hd7 ;
            rom[17986] = 8'hea ;
            rom[17987] = 8'hf9 ;
            rom[17988] = 8'hfa ;
            rom[17989] = 8'hf0 ;
            rom[17990] = 8'hf8 ;
            rom[17991] = 8'hfe ;
            rom[17992] = 8'hc7 ;
            rom[17993] = 8'hf1 ;
            rom[17994] = 8'h02 ;
            rom[17995] = 8'hdd ;
            rom[17996] = 8'h14 ;
            rom[17997] = 8'h03 ;
            rom[17998] = 8'hea ;
            rom[17999] = 8'hec ;
            rom[18000] = 8'hed ;
            rom[18001] = 8'h0c ;
            rom[18002] = 8'h1d ;
            rom[18003] = 8'h0e ;
            rom[18004] = 8'h0e ;
            rom[18005] = 8'hfc ;
            rom[18006] = 8'h26 ;
            rom[18007] = 8'hf8 ;
            rom[18008] = 8'hec ;
            rom[18009] = 8'h09 ;
            rom[18010] = 8'h08 ;
            rom[18011] = 8'h0b ;
            rom[18012] = 8'h13 ;
            rom[18013] = 8'he1 ;
            rom[18014] = 8'hf9 ;
            rom[18015] = 8'hfe ;
            rom[18016] = 8'hd5 ;
            rom[18017] = 8'h06 ;
            rom[18018] = 8'hfc ;
            rom[18019] = 8'h11 ;
            rom[18020] = 8'hfc ;
            rom[18021] = 8'h00 ;
            rom[18022] = 8'h17 ;
            rom[18023] = 8'h02 ;
            rom[18024] = 8'hff ;
            rom[18025] = 8'h37 ;
            rom[18026] = 8'hf3 ;
            rom[18027] = 8'he4 ;
            rom[18028] = 8'hf7 ;
            rom[18029] = 8'h1c ;
            rom[18030] = 8'hd2 ;
            rom[18031] = 8'h1c ;
            rom[18032] = 8'h15 ;
            rom[18033] = 8'h08 ;
            rom[18034] = 8'h0d ;
            rom[18035] = 8'h0d ;
            rom[18036] = 8'he9 ;
            rom[18037] = 8'h03 ;
            rom[18038] = 8'he4 ;
            rom[18039] = 8'hff ;
            rom[18040] = 8'h1e ;
            rom[18041] = 8'h1f ;
            rom[18042] = 8'h00 ;
            rom[18043] = 8'h08 ;
            rom[18044] = 8'hf0 ;
            rom[18045] = 8'hfa ;
            rom[18046] = 8'h1a ;
            rom[18047] = 8'h0b ;
            rom[18048] = 8'h03 ;
            rom[18049] = 8'h08 ;
            rom[18050] = 8'hdf ;
            rom[18051] = 8'h15 ;
            rom[18052] = 8'h16 ;
            rom[18053] = 8'h1c ;
            rom[18054] = 8'h15 ;
            rom[18055] = 8'h0e ;
            rom[18056] = 8'h24 ;
            rom[18057] = 8'he7 ;
            rom[18058] = 8'hea ;
            rom[18059] = 8'hee ;
            rom[18060] = 8'hf8 ;
            rom[18061] = 8'h16 ;
            rom[18062] = 8'h01 ;
            rom[18063] = 8'h1b ;
            rom[18064] = 8'h15 ;
            rom[18065] = 8'h2a ;
            rom[18066] = 8'hea ;
            rom[18067] = 8'hfb ;
            rom[18068] = 8'hf6 ;
            rom[18069] = 8'hfb ;
            rom[18070] = 8'hef ;
            rom[18071] = 8'h19 ;
            rom[18072] = 8'hfa ;
            rom[18073] = 8'hfe ;
            rom[18074] = 8'hf5 ;
            rom[18075] = 8'hed ;
            rom[18076] = 8'h06 ;
            rom[18077] = 8'hd0 ;
            rom[18078] = 8'hf5 ;
            rom[18079] = 8'hed ;
            rom[18080] = 8'hf9 ;
            rom[18081] = 8'he7 ;
            rom[18082] = 8'h0a ;
            rom[18083] = 8'hdd ;
            rom[18084] = 8'hce ;
            rom[18085] = 8'h20 ;
            rom[18086] = 8'hf9 ;
            rom[18087] = 8'h1d ;
            rom[18088] = 8'h0d ;
            rom[18089] = 8'he6 ;
            rom[18090] = 8'he8 ;
            rom[18091] = 8'hff ;
            rom[18092] = 8'h28 ;
            rom[18093] = 8'hd8 ;
            rom[18094] = 8'hef ;
            rom[18095] = 8'hed ;
            rom[18096] = 8'hf1 ;
            rom[18097] = 8'hdf ;
            rom[18098] = 8'hf9 ;
            rom[18099] = 8'hc6 ;
            rom[18100] = 8'hf1 ;
            rom[18101] = 8'h1b ;
            rom[18102] = 8'h3c ;
            rom[18103] = 8'hf5 ;
            rom[18104] = 8'h1a ;
            rom[18105] = 8'hcf ;
            rom[18106] = 8'h09 ;
            rom[18107] = 8'he8 ;
            rom[18108] = 8'h03 ;
            rom[18109] = 8'hf4 ;
            rom[18110] = 8'h14 ;
            rom[18111] = 8'hf0 ;
            rom[18112] = 8'h29 ;
            rom[18113] = 8'hb5 ;
            rom[18114] = 8'hf8 ;
            rom[18115] = 8'h0b ;
            rom[18116] = 8'h03 ;
            rom[18117] = 8'hee ;
            rom[18118] = 8'he4 ;
            rom[18119] = 8'he8 ;
            rom[18120] = 8'h20 ;
            rom[18121] = 8'hfc ;
            rom[18122] = 8'h08 ;
            rom[18123] = 8'hff ;
            rom[18124] = 8'h23 ;
            rom[18125] = 8'hd3 ;
            rom[18126] = 8'h0b ;
            rom[18127] = 8'h04 ;
            rom[18128] = 8'h09 ;
            rom[18129] = 8'h16 ;
            rom[18130] = 8'h0d ;
            rom[18131] = 8'h2e ;
            rom[18132] = 8'h10 ;
            rom[18133] = 8'hea ;
            rom[18134] = 8'hfd ;
            rom[18135] = 8'hd9 ;
            rom[18136] = 8'h24 ;
            rom[18137] = 8'he0 ;
            rom[18138] = 8'hdd ;
            rom[18139] = 8'hf2 ;
            rom[18140] = 8'he3 ;
            rom[18141] = 8'h2b ;
            rom[18142] = 8'hee ;
            rom[18143] = 8'h19 ;
            rom[18144] = 8'hf6 ;
            rom[18145] = 8'heb ;
            rom[18146] = 8'hf9 ;
            rom[18147] = 8'h06 ;
            rom[18148] = 8'hf4 ;
            rom[18149] = 8'hc6 ;
            rom[18150] = 8'hfd ;
            rom[18151] = 8'hc5 ;
            rom[18152] = 8'h25 ;
            rom[18153] = 8'h19 ;
            rom[18154] = 8'hec ;
            rom[18155] = 8'hfd ;
            rom[18156] = 8'hda ;
            rom[18157] = 8'hf2 ;
            rom[18158] = 8'hed ;
            rom[18159] = 8'hfd ;
            rom[18160] = 8'h35 ;
            rom[18161] = 8'hdf ;
            rom[18162] = 8'hf7 ;
            rom[18163] = 8'h09 ;
            rom[18164] = 8'h1b ;
            rom[18165] = 8'hf3 ;
            rom[18166] = 8'hfc ;
            rom[18167] = 8'h2d ;
            rom[18168] = 8'hd3 ;
            rom[18169] = 8'h22 ;
            rom[18170] = 8'h37 ;
            rom[18171] = 8'hef ;
            rom[18172] = 8'hee ;
            rom[18173] = 8'h0c ;
            rom[18174] = 8'he7 ;
            rom[18175] = 8'h07 ;
            rom[18176] = 8'hf6 ;
            rom[18177] = 8'hd8 ;
            rom[18178] = 8'hdd ;
            rom[18179] = 8'h26 ;
            rom[18180] = 8'hff ;
            rom[18181] = 8'hec ;
            rom[18182] = 8'h26 ;
            rom[18183] = 8'he9 ;
            rom[18184] = 8'h22 ;
            rom[18185] = 8'hd5 ;
            rom[18186] = 8'hff ;
            rom[18187] = 8'hc4 ;
            rom[18188] = 8'hed ;
            rom[18189] = 8'h01 ;
            rom[18190] = 8'hf9 ;
            rom[18191] = 8'hed ;
            rom[18192] = 8'he4 ;
            rom[18193] = 8'h15 ;
            rom[18194] = 8'h08 ;
            rom[18195] = 8'he9 ;
            rom[18196] = 8'h03 ;
            rom[18197] = 8'hed ;
            rom[18198] = 8'hf5 ;
            rom[18199] = 8'he5 ;
            rom[18200] = 8'hfe ;
            rom[18201] = 8'h06 ;
            rom[18202] = 8'h0c ;
            rom[18203] = 8'h02 ;
            rom[18204] = 8'h0b ;
            rom[18205] = 8'he6 ;
            rom[18206] = 8'h16 ;
            rom[18207] = 8'hc5 ;
            rom[18208] = 8'hf1 ;
            rom[18209] = 8'hfb ;
            rom[18210] = 8'hdd ;
            rom[18211] = 8'h0b ;
            rom[18212] = 8'hd1 ;
            rom[18213] = 8'h2a ;
            rom[18214] = 8'h00 ;
            rom[18215] = 8'h0b ;
            rom[18216] = 8'hda ;
            rom[18217] = 8'hd8 ;
            rom[18218] = 8'h08 ;
            rom[18219] = 8'hda ;
            rom[18220] = 8'h2b ;
            rom[18221] = 8'hf8 ;
            rom[18222] = 8'hf1 ;
            rom[18223] = 8'hf3 ;
            rom[18224] = 8'h17 ;
            rom[18225] = 8'hde ;
            rom[18226] = 8'h18 ;
            rom[18227] = 8'hbc ;
            rom[18228] = 8'h34 ;
            rom[18229] = 8'hf7 ;
            rom[18230] = 8'hda ;
            rom[18231] = 8'h17 ;
            rom[18232] = 8'h08 ;
            rom[18233] = 8'h05 ;
            rom[18234] = 8'h0b ;
            rom[18235] = 8'hd8 ;
            rom[18236] = 8'hf8 ;
            rom[18237] = 8'h19 ;
            rom[18238] = 8'he7 ;
            rom[18239] = 8'hcb ;
            rom[18240] = 8'hd3 ;
            rom[18241] = 8'hd6 ;
            rom[18242] = 8'hed ;
            rom[18243] = 8'h12 ;
            rom[18244] = 8'h10 ;
            rom[18245] = 8'h0a ;
            rom[18246] = 8'he3 ;
            rom[18247] = 8'hf4 ;
            rom[18248] = 8'h13 ;
            rom[18249] = 8'hde ;
            rom[18250] = 8'hfb ;
            rom[18251] = 8'h14 ;
            rom[18252] = 8'h29 ;
            rom[18253] = 8'hd2 ;
            rom[18254] = 8'h13 ;
            rom[18255] = 8'h0b ;
            rom[18256] = 8'h04 ;
            rom[18257] = 8'hed ;
            rom[18258] = 8'h10 ;
            rom[18259] = 8'he5 ;
            rom[18260] = 8'hfa ;
            rom[18261] = 8'hec ;
            rom[18262] = 8'hd8 ;
            rom[18263] = 8'h0c ;
            rom[18264] = 8'h22 ;
            rom[18265] = 8'hf6 ;
            rom[18266] = 8'h10 ;
            rom[18267] = 8'h03 ;
            rom[18268] = 8'hff ;
            rom[18269] = 8'h09 ;
            rom[18270] = 8'hea ;
            rom[18271] = 8'h0f ;
            rom[18272] = 8'hdd ;
            rom[18273] = 8'hde ;
            rom[18274] = 8'hf2 ;
            rom[18275] = 8'h2a ;
            rom[18276] = 8'h0e ;
            rom[18277] = 8'h02 ;
            rom[18278] = 8'h12 ;
            rom[18279] = 8'hef ;
            rom[18280] = 8'he9 ;
            rom[18281] = 8'he3 ;
            rom[18282] = 8'hf6 ;
            rom[18283] = 8'h1a ;
            rom[18284] = 8'hf3 ;
            rom[18285] = 8'h09 ;
            rom[18286] = 8'hf6 ;
            rom[18287] = 8'hfb ;
            rom[18288] = 8'hf5 ;
            rom[18289] = 8'he9 ;
            rom[18290] = 8'h0e ;
            rom[18291] = 8'hd0 ;
            rom[18292] = 8'hff ;
            rom[18293] = 8'h07 ;
            rom[18294] = 8'h0a ;
            rom[18295] = 8'h2a ;
            rom[18296] = 8'hd9 ;
            rom[18297] = 8'h01 ;
            rom[18298] = 8'h0c ;
            rom[18299] = 8'h1f ;
            rom[18300] = 8'hdd ;
            rom[18301] = 8'h0f ;
            rom[18302] = 8'he1 ;
            rom[18303] = 8'hfa ;
            rom[18304] = 8'hd6 ;
            rom[18305] = 8'he5 ;
            rom[18306] = 8'hf4 ;
            rom[18307] = 8'h1c ;
            rom[18308] = 8'h03 ;
            rom[18309] = 8'h03 ;
            rom[18310] = 8'h0e ;
            rom[18311] = 8'hfb ;
            rom[18312] = 8'hd5 ;
            rom[18313] = 8'hdd ;
            rom[18314] = 8'h1d ;
            rom[18315] = 8'hf2 ;
            rom[18316] = 8'hf5 ;
            rom[18317] = 8'hf6 ;
            rom[18318] = 8'hf4 ;
            rom[18319] = 8'h0b ;
            rom[18320] = 8'h06 ;
            rom[18321] = 8'h08 ;
            rom[18322] = 8'h10 ;
            rom[18323] = 8'hdc ;
            rom[18324] = 8'h13 ;
            rom[18325] = 8'hfb ;
            rom[18326] = 8'hdc ;
            rom[18327] = 8'h0d ;
            rom[18328] = 8'h2a ;
            rom[18329] = 8'h08 ;
            rom[18330] = 8'h25 ;
            rom[18331] = 8'hee ;
            rom[18332] = 8'hfe ;
            rom[18333] = 8'hf8 ;
            rom[18334] = 8'h17 ;
            rom[18335] = 8'h13 ;
            rom[18336] = 8'h1f ;
            rom[18337] = 8'hf9 ;
            rom[18338] = 8'h30 ;
            rom[18339] = 8'h02 ;
            rom[18340] = 8'h0e ;
            rom[18341] = 8'h20 ;
            rom[18342] = 8'hf3 ;
            rom[18343] = 8'he4 ;
            rom[18344] = 8'h00 ;
            rom[18345] = 8'h01 ;
            rom[18346] = 8'hf7 ;
            rom[18347] = 8'h11 ;
            rom[18348] = 8'h06 ;
            rom[18349] = 8'h18 ;
            rom[18350] = 8'hd9 ;
            rom[18351] = 8'hf6 ;
            rom[18352] = 8'h08 ;
            rom[18353] = 8'h1a ;
            rom[18354] = 8'he4 ;
            rom[18355] = 8'h09 ;
            rom[18356] = 8'he5 ;
            rom[18357] = 8'hfd ;
            rom[18358] = 8'hfa ;
            rom[18359] = 8'hf1 ;
            rom[18360] = 8'h16 ;
            rom[18361] = 8'hef ;
            rom[18362] = 8'h02 ;
            rom[18363] = 8'he4 ;
            rom[18364] = 8'h07 ;
            rom[18365] = 8'hf0 ;
            rom[18366] = 8'h08 ;
            rom[18367] = 8'h06 ;
            rom[18368] = 8'hda ;
            rom[18369] = 8'hf0 ;
            rom[18370] = 8'h07 ;
            rom[18371] = 8'h04 ;
            rom[18372] = 8'hfe ;
            rom[18373] = 8'hfe ;
            rom[18374] = 8'hef ;
            rom[18375] = 8'h17 ;
            rom[18376] = 8'hf1 ;
            rom[18377] = 8'he3 ;
            rom[18378] = 8'h05 ;
            rom[18379] = 8'hfe ;
            rom[18380] = 8'h1a ;
            rom[18381] = 8'hde ;
            rom[18382] = 8'h04 ;
            rom[18383] = 8'hf4 ;
            rom[18384] = 8'h2f ;
            rom[18385] = 8'hfc ;
            rom[18386] = 8'hed ;
            rom[18387] = 8'h24 ;
            rom[18388] = 8'hd1 ;
            rom[18389] = 8'hf5 ;
            rom[18390] = 8'h18 ;
            rom[18391] = 8'hf1 ;
            rom[18392] = 8'h0a ;
            rom[18393] = 8'hf8 ;
            rom[18394] = 8'h04 ;
            rom[18395] = 8'h20 ;
            rom[18396] = 8'he6 ;
            rom[18397] = 8'h32 ;
            rom[18398] = 8'hfe ;
            rom[18399] = 8'hfc ;
            rom[18400] = 8'h19 ;
            rom[18401] = 8'h1d ;
            rom[18402] = 8'he5 ;
            rom[18403] = 8'h07 ;
            rom[18404] = 8'hf5 ;
            rom[18405] = 8'h3e ;
            rom[18406] = 8'h39 ;
            rom[18407] = 8'hee ;
            rom[18408] = 8'hff ;
            rom[18409] = 8'hf3 ;
            rom[18410] = 8'h12 ;
            rom[18411] = 8'h05 ;
            rom[18412] = 8'hee ;
            rom[18413] = 8'hc3 ;
            rom[18414] = 8'hd7 ;
            rom[18415] = 8'hfd ;
            rom[18416] = 8'h0f ;
            rom[18417] = 8'hea ;
            rom[18418] = 8'h11 ;
            rom[18419] = 8'h01 ;
            rom[18420] = 8'he0 ;
            rom[18421] = 8'hfe ;
            rom[18422] = 8'hf4 ;
            rom[18423] = 8'hf4 ;
            rom[18424] = 8'he9 ;
            rom[18425] = 8'h13 ;
            rom[18426] = 8'hfb ;
            rom[18427] = 8'he3 ;
            rom[18428] = 8'h1b ;
            rom[18429] = 8'h1e ;
            rom[18430] = 8'hfc ;
            rom[18431] = 8'h1b ;
            rom[18432] = 8'h02 ;
            rom[18433] = 8'hf3 ;
            rom[18434] = 8'hfa ;
            rom[18435] = 8'h0d ;
            rom[18436] = 8'hd7 ;
            rom[18437] = 8'h23 ;
            rom[18438] = 8'h09 ;
            rom[18439] = 8'h03 ;
            rom[18440] = 8'h1e ;
            rom[18441] = 8'hdd ;
            rom[18442] = 8'hd2 ;
            rom[18443] = 8'hf9 ;
            rom[18444] = 8'hfb ;
            rom[18445] = 8'hd8 ;
            rom[18446] = 8'hd2 ;
            rom[18447] = 8'h1c ;
            rom[18448] = 8'hf2 ;
            rom[18449] = 8'h16 ;
            rom[18450] = 8'h0c ;
            rom[18451] = 8'h0c ;
            rom[18452] = 8'h0a ;
            rom[18453] = 8'h13 ;
            rom[18454] = 8'hcc ;
            rom[18455] = 8'h15 ;
            rom[18456] = 8'hf8 ;
            rom[18457] = 8'hf0 ;
            rom[18458] = 8'h01 ;
            rom[18459] = 8'hff ;
            rom[18460] = 8'hf5 ;
            rom[18461] = 8'h0b ;
            rom[18462] = 8'h15 ;
            rom[18463] = 8'he9 ;
            rom[18464] = 8'h0f ;
            rom[18465] = 8'hf8 ;
            rom[18466] = 8'h0b ;
            rom[18467] = 8'hf6 ;
            rom[18468] = 8'hc9 ;
            rom[18469] = 8'h18 ;
            rom[18470] = 8'h08 ;
            rom[18471] = 8'hf7 ;
            rom[18472] = 8'h05 ;
            rom[18473] = 8'hd7 ;
            rom[18474] = 8'h0a ;
            rom[18475] = 8'h03 ;
            rom[18476] = 8'hf5 ;
            rom[18477] = 8'hcc ;
            rom[18478] = 8'hf4 ;
            rom[18479] = 8'h20 ;
            rom[18480] = 8'hf3 ;
            rom[18481] = 8'hfa ;
            rom[18482] = 8'h09 ;
            rom[18483] = 8'h12 ;
            rom[18484] = 8'h14 ;
            rom[18485] = 8'h1b ;
            rom[18486] = 8'h23 ;
            rom[18487] = 8'h01 ;
            rom[18488] = 8'he7 ;
            rom[18489] = 8'hf4 ;
            rom[18490] = 8'h19 ;
            rom[18491] = 8'hdf ;
            rom[18492] = 8'hf1 ;
            rom[18493] = 8'hf9 ;
            rom[18494] = 8'h16 ;
            rom[18495] = 8'h0d ;
            rom[18496] = 8'h23 ;
            rom[18497] = 8'h08 ;
            rom[18498] = 8'h0c ;
            rom[18499] = 8'hf4 ;
            rom[18500] = 8'he4 ;
            rom[18501] = 8'hf3 ;
            rom[18502] = 8'hf7 ;
            rom[18503] = 8'hd3 ;
            rom[18504] = 8'hf0 ;
            rom[18505] = 8'h0e ;
            rom[18506] = 8'hcb ;
            rom[18507] = 8'hcd ;
            rom[18508] = 8'h13 ;
            rom[18509] = 8'he7 ;
            rom[18510] = 8'h0a ;
            rom[18511] = 8'h2a ;
            rom[18512] = 8'h1a ;
            rom[18513] = 8'he1 ;
            rom[18514] = 8'hf1 ;
            rom[18515] = 8'hf6 ;
            rom[18516] = 8'hbf ;
            rom[18517] = 8'hed ;
            rom[18518] = 8'h1c ;
            rom[18519] = 8'h36 ;
            rom[18520] = 8'h1b ;
            rom[18521] = 8'h0e ;
            rom[18522] = 8'h18 ;
            rom[18523] = 8'heb ;
            rom[18524] = 8'h09 ;
            rom[18525] = 8'hf4 ;
            rom[18526] = 8'h0c ;
            rom[18527] = 8'h02 ;
            rom[18528] = 8'h26 ;
            rom[18529] = 8'hff ;
            rom[18530] = 8'h00 ;
            rom[18531] = 8'heb ;
            rom[18532] = 8'he2 ;
            rom[18533] = 8'he8 ;
            rom[18534] = 8'hf6 ;
            rom[18535] = 8'h0c ;
            rom[18536] = 8'h2a ;
            rom[18537] = 8'hef ;
            rom[18538] = 8'h20 ;
            rom[18539] = 8'h00 ;
            rom[18540] = 8'hf2 ;
            rom[18541] = 8'he6 ;
            rom[18542] = 8'hf2 ;
            rom[18543] = 8'h0c ;
            rom[18544] = 8'h08 ;
            rom[18545] = 8'hea ;
            rom[18546] = 8'hed ;
            rom[18547] = 8'h0d ;
            rom[18548] = 8'h15 ;
            rom[18549] = 8'h0b ;
            rom[18550] = 8'hda ;
            rom[18551] = 8'h14 ;
            rom[18552] = 8'h0d ;
            rom[18553] = 8'h0e ;
            rom[18554] = 8'hf4 ;
            rom[18555] = 8'he2 ;
            rom[18556] = 8'hfb ;
            rom[18557] = 8'h18 ;
            rom[18558] = 8'h0a ;
            rom[18559] = 8'h0b ;
            rom[18560] = 8'h11 ;
            rom[18561] = 8'hf2 ;
            rom[18562] = 8'h04 ;
            rom[18563] = 8'hfd ;
            rom[18564] = 8'h0a ;
            rom[18565] = 8'h0d ;
            rom[18566] = 8'h07 ;
            rom[18567] = 8'h23 ;
            rom[18568] = 8'hf5 ;
            rom[18569] = 8'hfe ;
            rom[18570] = 8'h0b ;
            rom[18571] = 8'h14 ;
            rom[18572] = 8'h02 ;
            rom[18573] = 8'h02 ;
            rom[18574] = 8'h11 ;
            rom[18575] = 8'h05 ;
            rom[18576] = 8'h03 ;
            rom[18577] = 8'h00 ;
            rom[18578] = 8'h13 ;
            rom[18579] = 8'h09 ;
            rom[18580] = 8'h10 ;
            rom[18581] = 8'h0a ;
            rom[18582] = 8'h22 ;
            rom[18583] = 8'hcd ;
            rom[18584] = 8'h11 ;
            rom[18585] = 8'h17 ;
            rom[18586] = 8'hf9 ;
            rom[18587] = 8'heb ;
            rom[18588] = 8'he3 ;
            rom[18589] = 8'h00 ;
            rom[18590] = 8'h06 ;
            rom[18591] = 8'h0c ;
            rom[18592] = 8'he9 ;
            rom[18593] = 8'hfe ;
            rom[18594] = 8'hf5 ;
            rom[18595] = 8'hcf ;
            rom[18596] = 8'hdf ;
            rom[18597] = 8'h29 ;
            rom[18598] = 8'h10 ;
            rom[18599] = 8'he1 ;
            rom[18600] = 8'he4 ;
            rom[18601] = 8'hc9 ;
            rom[18602] = 8'h0a ;
            rom[18603] = 8'hec ;
            rom[18604] = 8'h02 ;
            rom[18605] = 8'h0c ;
            rom[18606] = 8'h23 ;
            rom[18607] = 8'hf3 ;
            rom[18608] = 8'hfa ;
            rom[18609] = 8'hd8 ;
            rom[18610] = 8'h11 ;
            rom[18611] = 8'he6 ;
            rom[18612] = 8'he6 ;
            rom[18613] = 8'h0a ;
            rom[18614] = 8'h0a ;
            rom[18615] = 8'h0c ;
            rom[18616] = 8'hef ;
            rom[18617] = 8'he4 ;
            rom[18618] = 8'h0f ;
            rom[18619] = 8'he0 ;
            rom[18620] = 8'hf9 ;
            rom[18621] = 8'he3 ;
            rom[18622] = 8'h09 ;
            rom[18623] = 8'h10 ;
            rom[18624] = 8'h01 ;
            rom[18625] = 8'hf8 ;
            rom[18626] = 8'hd0 ;
            rom[18627] = 8'he2 ;
            rom[18628] = 8'h03 ;
            rom[18629] = 8'hfe ;
            rom[18630] = 8'hea ;
            rom[18631] = 8'h0e ;
            rom[18632] = 8'hf3 ;
            rom[18633] = 8'hdf ;
            rom[18634] = 8'hd6 ;
            rom[18635] = 8'h11 ;
            rom[18636] = 8'hce ;
            rom[18637] = 8'hfd ;
            rom[18638] = 8'hf4 ;
            rom[18639] = 8'h13 ;
            rom[18640] = 8'hf5 ;
            rom[18641] = 8'h1f ;
            rom[18642] = 8'h0c ;
            rom[18643] = 8'hed ;
            rom[18644] = 8'heb ;
            rom[18645] = 8'h23 ;
            rom[18646] = 8'h07 ;
            rom[18647] = 8'h17 ;
            rom[18648] = 8'hf3 ;
            rom[18649] = 8'h15 ;
            rom[18650] = 8'h0e ;
            rom[18651] = 8'h03 ;
            rom[18652] = 8'h14 ;
            rom[18653] = 8'hed ;
            rom[18654] = 8'h12 ;
            rom[18655] = 8'h04 ;
            rom[18656] = 8'he5 ;
            rom[18657] = 8'h0c ;
            rom[18658] = 8'h08 ;
            rom[18659] = 8'h23 ;
            rom[18660] = 8'hed ;
            rom[18661] = 8'h04 ;
            rom[18662] = 8'hf9 ;
            rom[18663] = 8'h00 ;
            rom[18664] = 8'hfb ;
            rom[18665] = 8'h0a ;
            rom[18666] = 8'hf9 ;
            rom[18667] = 8'heb ;
            rom[18668] = 8'h0c ;
            rom[18669] = 8'hfc ;
            rom[18670] = 8'h12 ;
            rom[18671] = 8'h0a ;
            rom[18672] = 8'h06 ;
            rom[18673] = 8'hfd ;
            rom[18674] = 8'he8 ;
            rom[18675] = 8'h0e ;
            rom[18676] = 8'hf0 ;
            rom[18677] = 8'hf5 ;
            rom[18678] = 8'h08 ;
            rom[18679] = 8'h04 ;
            rom[18680] = 8'h16 ;
            rom[18681] = 8'hfe ;
            rom[18682] = 8'he8 ;
            rom[18683] = 8'h15 ;
            rom[18684] = 8'h08 ;
            rom[18685] = 8'h06 ;
            rom[18686] = 8'hff ;
            rom[18687] = 8'h32 ;
            rom[18688] = 8'hed ;
            rom[18689] = 8'hea ;
            rom[18690] = 8'hf1 ;
            rom[18691] = 8'he6 ;
            rom[18692] = 8'h12 ;
            rom[18693] = 8'h05 ;
            rom[18694] = 8'hee ;
            rom[18695] = 8'hdd ;
            rom[18696] = 8'h00 ;
            rom[18697] = 8'hf3 ;
            rom[18698] = 8'h2b ;
            rom[18699] = 8'h19 ;
            rom[18700] = 8'h01 ;
            rom[18701] = 8'h0e ;
            rom[18702] = 8'hf4 ;
            rom[18703] = 8'h07 ;
            rom[18704] = 8'h05 ;
            rom[18705] = 8'h19 ;
            rom[18706] = 8'hfa ;
            rom[18707] = 8'h05 ;
            rom[18708] = 8'h10 ;
            rom[18709] = 8'heb ;
            rom[18710] = 8'hfa ;
            rom[18711] = 8'hf3 ;
            rom[18712] = 8'hf1 ;
            rom[18713] = 8'h0a ;
            rom[18714] = 8'hd4 ;
            rom[18715] = 8'he9 ;
            rom[18716] = 8'he5 ;
            rom[18717] = 8'hf8 ;
            rom[18718] = 8'h1c ;
            rom[18719] = 8'hd4 ;
            rom[18720] = 8'h0e ;
            rom[18721] = 8'hf9 ;
            rom[18722] = 8'hdb ;
            rom[18723] = 8'hfe ;
            rom[18724] = 8'hf0 ;
            rom[18725] = 8'h2f ;
            rom[18726] = 8'hf6 ;
            rom[18727] = 8'h01 ;
            rom[18728] = 8'hec ;
            rom[18729] = 8'hf2 ;
            rom[18730] = 8'hf4 ;
            rom[18731] = 8'hfd ;
            rom[18732] = 8'hee ;
            rom[18733] = 8'hfb ;
            rom[18734] = 8'h17 ;
            rom[18735] = 8'he8 ;
            rom[18736] = 8'h1b ;
            rom[18737] = 8'hd2 ;
            rom[18738] = 8'he2 ;
            rom[18739] = 8'h22 ;
            rom[18740] = 8'hf4 ;
            rom[18741] = 8'h0b ;
            rom[18742] = 8'hd7 ;
            rom[18743] = 8'he1 ;
            rom[18744] = 8'hd9 ;
            rom[18745] = 8'heb ;
            rom[18746] = 8'he7 ;
            rom[18747] = 8'h26 ;
            rom[18748] = 8'h0e ;
            rom[18749] = 8'h06 ;
            rom[18750] = 8'h03 ;
            rom[18751] = 8'hfd ;
            rom[18752] = 8'hff ;
            rom[18753] = 8'h21 ;
            rom[18754] = 8'h0b ;
            rom[18755] = 8'hf5 ;
            rom[18756] = 8'he3 ;
            rom[18757] = 8'hf6 ;
            rom[18758] = 8'hfd ;
            rom[18759] = 8'h13 ;
            rom[18760] = 8'h11 ;
            rom[18761] = 8'hf2 ;
            rom[18762] = 8'he0 ;
            rom[18763] = 8'hfd ;
            rom[18764] = 8'h19 ;
            rom[18765] = 8'he7 ;
            rom[18766] = 8'h1a ;
            rom[18767] = 8'h08 ;
            rom[18768] = 8'h13 ;
            rom[18769] = 8'h12 ;
            rom[18770] = 8'h2e ;
            rom[18771] = 8'h23 ;
            rom[18772] = 8'hd7 ;
            rom[18773] = 8'hf9 ;
            rom[18774] = 8'h14 ;
            rom[18775] = 8'hfb ;
            rom[18776] = 8'h00 ;
            rom[18777] = 8'h19 ;
            rom[18778] = 8'hfd ;
            rom[18779] = 8'h0c ;
            rom[18780] = 8'hee ;
            rom[18781] = 8'h15 ;
            rom[18782] = 8'hf7 ;
            rom[18783] = 8'hfa ;
            rom[18784] = 8'h00 ;
            rom[18785] = 8'hfc ;
            rom[18786] = 8'heb ;
            rom[18787] = 8'hed ;
            rom[18788] = 8'hee ;
            rom[18789] = 8'h20 ;
            rom[18790] = 8'h09 ;
            rom[18791] = 8'hf6 ;
            rom[18792] = 8'hfb ;
            rom[18793] = 8'h0b ;
            rom[18794] = 8'h0e ;
            rom[18795] = 8'h11 ;
            rom[18796] = 8'h16 ;
            rom[18797] = 8'hdb ;
            rom[18798] = 8'h1e ;
            rom[18799] = 8'hfe ;
            rom[18800] = 8'hba ;
            rom[18801] = 8'h05 ;
            rom[18802] = 8'h0b ;
            rom[18803] = 8'h02 ;
            rom[18804] = 8'h05 ;
            rom[18805] = 8'h2c ;
            rom[18806] = 8'h06 ;
            rom[18807] = 8'h0c ;
            rom[18808] = 8'hf4 ;
            rom[18809] = 8'hfa ;
            rom[18810] = 8'hf8 ;
            rom[18811] = 8'hff ;
            rom[18812] = 8'he0 ;
            rom[18813] = 8'h14 ;
            rom[18814] = 8'h12 ;
            rom[18815] = 8'hf4 ;
            rom[18816] = 8'hfb ;
            rom[18817] = 8'hfb ;
            rom[18818] = 8'hf9 ;
            rom[18819] = 8'h27 ;
            rom[18820] = 8'hd5 ;
            rom[18821] = 8'h06 ;
            rom[18822] = 8'h04 ;
            rom[18823] = 8'h09 ;
            rom[18824] = 8'h2c ;
            rom[18825] = 8'hee ;
            rom[18826] = 8'he2 ;
            rom[18827] = 8'hb4 ;
            rom[18828] = 8'h15 ;
            rom[18829] = 8'h0f ;
            rom[18830] = 8'h0d ;
            rom[18831] = 8'h1a ;
            rom[18832] = 8'hed ;
            rom[18833] = 8'h0d ;
            rom[18834] = 8'h16 ;
            rom[18835] = 8'hff ;
            rom[18836] = 8'h07 ;
            rom[18837] = 8'h11 ;
            rom[18838] = 8'hd9 ;
            rom[18839] = 8'h03 ;
            rom[18840] = 8'h05 ;
            rom[18841] = 8'h03 ;
            rom[18842] = 8'h14 ;
            rom[18843] = 8'h0e ;
            rom[18844] = 8'he9 ;
            rom[18845] = 8'hf8 ;
            rom[18846] = 8'h05 ;
            rom[18847] = 8'he7 ;
            rom[18848] = 8'he3 ;
            rom[18849] = 8'hf8 ;
            rom[18850] = 8'hf9 ;
            rom[18851] = 8'h04 ;
            rom[18852] = 8'hcd ;
            rom[18853] = 8'h06 ;
            rom[18854] = 8'h10 ;
            rom[18855] = 8'he5 ;
            rom[18856] = 8'h09 ;
            rom[18857] = 8'h13 ;
            rom[18858] = 8'h27 ;
            rom[18859] = 8'h06 ;
            rom[18860] = 8'hdf ;
            rom[18861] = 8'hde ;
            rom[18862] = 8'hd3 ;
            rom[18863] = 8'h1f ;
            rom[18864] = 8'hd6 ;
            rom[18865] = 8'h10 ;
            rom[18866] = 8'h21 ;
            rom[18867] = 8'h09 ;
            rom[18868] = 8'h0f ;
            rom[18869] = 8'h07 ;
            rom[18870] = 8'hf5 ;
            rom[18871] = 8'hf5 ;
            rom[18872] = 8'hfe ;
            rom[18873] = 8'he5 ;
            rom[18874] = 8'hfd ;
            rom[18875] = 8'hc3 ;
            rom[18876] = 8'h0f ;
            rom[18877] = 8'h03 ;
            rom[18878] = 8'hda ;
            rom[18879] = 8'h04 ;
            rom[18880] = 8'hfa ;
            rom[18881] = 8'h01 ;
            rom[18882] = 8'h12 ;
            rom[18883] = 8'hfa ;
            rom[18884] = 8'h0a ;
            rom[18885] = 8'hfe ;
            rom[18886] = 8'hed ;
            rom[18887] = 8'hdc ;
            rom[18888] = 8'h31 ;
            rom[18889] = 8'h0e ;
            rom[18890] = 8'hcc ;
            rom[18891] = 8'hf9 ;
            rom[18892] = 8'h26 ;
            rom[18893] = 8'h18 ;
            rom[18894] = 8'hfd ;
            rom[18895] = 8'h03 ;
            rom[18896] = 8'h03 ;
            rom[18897] = 8'h13 ;
            rom[18898] = 8'hf5 ;
            rom[18899] = 8'h21 ;
            rom[18900] = 8'hd6 ;
            rom[18901] = 8'h02 ;
            rom[18902] = 8'hfe ;
            rom[18903] = 8'hff ;
            rom[18904] = 8'h1e ;
            rom[18905] = 8'hf0 ;
            rom[18906] = 8'he4 ;
            rom[18907] = 8'hff ;
            rom[18908] = 8'h10 ;
            rom[18909] = 8'hee ;
            rom[18910] = 8'h0a ;
            rom[18911] = 8'hed ;
            rom[18912] = 8'h13 ;
            rom[18913] = 8'h14 ;
            rom[18914] = 8'hf4 ;
            rom[18915] = 8'h08 ;
            rom[18916] = 8'hde ;
            rom[18917] = 8'h0d ;
            rom[18918] = 8'h1f ;
            rom[18919] = 8'h18 ;
            rom[18920] = 8'h13 ;
            rom[18921] = 8'h11 ;
            rom[18922] = 8'h1f ;
            rom[18923] = 8'hec ;
            rom[18924] = 8'hf9 ;
            rom[18925] = 8'h03 ;
            rom[18926] = 8'h00 ;
            rom[18927] = 8'he0 ;
            rom[18928] = 8'he6 ;
            rom[18929] = 8'hce ;
            rom[18930] = 8'hde ;
            rom[18931] = 8'he6 ;
            rom[18932] = 8'h0a ;
            rom[18933] = 8'heb ;
            rom[18934] = 8'hfb ;
            rom[18935] = 8'hf7 ;
            rom[18936] = 8'hbb ;
            rom[18937] = 8'hf0 ;
            rom[18938] = 8'h23 ;
            rom[18939] = 8'h1c ;
            rom[18940] = 8'hfc ;
            rom[18941] = 8'he9 ;
            rom[18942] = 8'hf9 ;
            rom[18943] = 8'hf6 ;
            rom[18944] = 8'h02 ;
            rom[18945] = 8'he7 ;
            rom[18946] = 8'hff ;
            rom[18947] = 8'hff ;
            rom[18948] = 8'hfd ;
            rom[18949] = 8'hc2 ;
            rom[18950] = 8'h10 ;
            rom[18951] = 8'hde ;
            rom[18952] = 8'h0b ;
            rom[18953] = 8'h05 ;
            rom[18954] = 8'hf6 ;
            rom[18955] = 8'hd8 ;
            rom[18956] = 8'hd3 ;
            rom[18957] = 8'hec ;
            rom[18958] = 8'hd1 ;
            rom[18959] = 8'hd5 ;
            rom[18960] = 8'he9 ;
            rom[18961] = 8'h00 ;
            rom[18962] = 8'hc6 ;
            rom[18963] = 8'hd6 ;
            rom[18964] = 8'h24 ;
            rom[18965] = 8'he9 ;
            rom[18966] = 8'hf5 ;
            rom[18967] = 8'hbc ;
            rom[18968] = 8'h0f ;
            rom[18969] = 8'h0d ;
            rom[18970] = 8'h02 ;
            rom[18971] = 8'hee ;
            rom[18972] = 8'h13 ;
            rom[18973] = 8'h1a ;
            rom[18974] = 8'h06 ;
            rom[18975] = 8'hfe ;
            rom[18976] = 8'h05 ;
            rom[18977] = 8'h0d ;
            rom[18978] = 8'hfa ;
            rom[18979] = 8'he9 ;
            rom[18980] = 8'h2a ;
            rom[18981] = 8'he6 ;
            rom[18982] = 8'hcd ;
            rom[18983] = 8'h0a ;
            rom[18984] = 8'h01 ;
            rom[18985] = 8'h10 ;
            rom[18986] = 8'hea ;
            rom[18987] = 8'hc3 ;
            rom[18988] = 8'h06 ;
            rom[18989] = 8'h08 ;
            rom[18990] = 8'h00 ;
            rom[18991] = 8'hdc ;
            rom[18992] = 8'hd9 ;
            rom[18993] = 8'h15 ;
            rom[18994] = 8'hda ;
            rom[18995] = 8'he7 ;
            rom[18996] = 8'h06 ;
            rom[18997] = 8'h14 ;
            rom[18998] = 8'he8 ;
            rom[18999] = 8'h09 ;
            rom[19000] = 8'h1a ;
            rom[19001] = 8'h12 ;
            rom[19002] = 8'h06 ;
            rom[19003] = 8'h09 ;
            rom[19004] = 8'hef ;
            rom[19005] = 8'hfe ;
            rom[19006] = 8'hd7 ;
            rom[19007] = 8'hdb ;
            rom[19008] = 8'h19 ;
            rom[19009] = 8'he0 ;
            rom[19010] = 8'h23 ;
            rom[19011] = 8'hff ;
            rom[19012] = 8'h23 ;
            rom[19013] = 8'h0d ;
            rom[19014] = 8'he8 ;
            rom[19015] = 8'h09 ;
            rom[19016] = 8'h21 ;
            rom[19017] = 8'hfa ;
            rom[19018] = 8'hf3 ;
            rom[19019] = 8'h21 ;
            rom[19020] = 8'h01 ;
            rom[19021] = 8'hd0 ;
            rom[19022] = 8'hf4 ;
            rom[19023] = 8'h02 ;
            rom[19024] = 8'hdf ;
            rom[19025] = 8'hdd ;
            rom[19026] = 8'hf5 ;
            rom[19027] = 8'hfa ;
            rom[19028] = 8'heb ;
            rom[19029] = 8'hf8 ;
            rom[19030] = 8'he3 ;
            rom[19031] = 8'h24 ;
            rom[19032] = 8'h04 ;
            rom[19033] = 8'hf5 ;
            rom[19034] = 8'h01 ;
            rom[19035] = 8'heb ;
            rom[19036] = 8'hf9 ;
            rom[19037] = 8'h11 ;
            rom[19038] = 8'h00 ;
            rom[19039] = 8'hf7 ;
            rom[19040] = 8'hff ;
            rom[19041] = 8'hb1 ;
            rom[19042] = 8'hf6 ;
            rom[19043] = 8'h08 ;
            rom[19044] = 8'hed ;
            rom[19045] = 8'hfd ;
            rom[19046] = 8'hdf ;
            rom[19047] = 8'hd1 ;
            rom[19048] = 8'hfe ;
            rom[19049] = 8'he2 ;
            rom[19050] = 8'hee ;
            rom[19051] = 8'h00 ;
            rom[19052] = 8'h16 ;
            rom[19053] = 8'h0b ;
            rom[19054] = 8'h07 ;
            rom[19055] = 8'hf9 ;
            rom[19056] = 8'hfc ;
            rom[19057] = 8'hf3 ;
            rom[19058] = 8'h08 ;
            rom[19059] = 8'hcc ;
            rom[19060] = 8'hfc ;
            rom[19061] = 8'hfc ;
            rom[19062] = 8'hfe ;
            rom[19063] = 8'hf3 ;
            rom[19064] = 8'hd4 ;
            rom[19065] = 8'hfd ;
            rom[19066] = 8'hf5 ;
            rom[19067] = 8'hd9 ;
            rom[19068] = 8'hde ;
            rom[19069] = 8'hcf ;
            rom[19070] = 8'hd0 ;
            rom[19071] = 8'hee ;
            rom[19072] = 8'hf4 ;
            rom[19073] = 8'h1c ;
            rom[19074] = 8'hfe ;
            rom[19075] = 8'hfc ;
            rom[19076] = 8'h05 ;
            rom[19077] = 8'he4 ;
            rom[19078] = 8'h21 ;
            rom[19079] = 8'h04 ;
            rom[19080] = 8'hfc ;
            rom[19081] = 8'h0d ;
            rom[19082] = 8'h11 ;
            rom[19083] = 8'h01 ;
            rom[19084] = 8'he9 ;
            rom[19085] = 8'h19 ;
            rom[19086] = 8'he7 ;
            rom[19087] = 8'h35 ;
            rom[19088] = 8'hf4 ;
            rom[19089] = 8'hd8 ;
            rom[19090] = 8'h0f ;
            rom[19091] = 8'hdd ;
            rom[19092] = 8'h0e ;
            rom[19093] = 8'h08 ;
            rom[19094] = 8'hf5 ;
            rom[19095] = 8'h15 ;
            rom[19096] = 8'he1 ;
            rom[19097] = 8'h11 ;
            rom[19098] = 8'h0c ;
            rom[19099] = 8'h0d ;
            rom[19100] = 8'h0e ;
            rom[19101] = 8'h16 ;
            rom[19102] = 8'h0b ;
            rom[19103] = 8'h19 ;
            rom[19104] = 8'h0b ;
            rom[19105] = 8'h01 ;
            rom[19106] = 8'hfc ;
            rom[19107] = 8'hb9 ;
            rom[19108] = 8'hf1 ;
            rom[19109] = 8'h00 ;
            rom[19110] = 8'hf9 ;
            rom[19111] = 8'h15 ;
            rom[19112] = 8'h2a ;
            rom[19113] = 8'hf5 ;
            rom[19114] = 8'hde ;
            rom[19115] = 8'h17 ;
            rom[19116] = 8'hf8 ;
            rom[19117] = 8'h05 ;
            rom[19118] = 8'h08 ;
            rom[19119] = 8'hef ;
            rom[19120] = 8'hf9 ;
            rom[19121] = 8'h04 ;
            rom[19122] = 8'hf5 ;
            rom[19123] = 8'h0c ;
            rom[19124] = 8'hfc ;
            rom[19125] = 8'he1 ;
            rom[19126] = 8'hf9 ;
            rom[19127] = 8'he5 ;
            rom[19128] = 8'h0f ;
            rom[19129] = 8'h1c ;
            rom[19130] = 8'h09 ;
            rom[19131] = 8'hd0 ;
            rom[19132] = 8'he4 ;
            rom[19133] = 8'h06 ;
            rom[19134] = 8'h17 ;
            rom[19135] = 8'h1b ;
            rom[19136] = 8'hd3 ;
            rom[19137] = 8'h08 ;
            rom[19138] = 8'hf7 ;
            rom[19139] = 8'h04 ;
            rom[19140] = 8'hd3 ;
            rom[19141] = 8'hf7 ;
            rom[19142] = 8'hd1 ;
            rom[19143] = 8'h23 ;
            rom[19144] = 8'hbc ;
            rom[19145] = 8'hdc ;
            rom[19146] = 8'h0c ;
            rom[19147] = 8'h2e ;
            rom[19148] = 8'hf0 ;
            rom[19149] = 8'hd6 ;
            rom[19150] = 8'he9 ;
            rom[19151] = 8'h08 ;
            rom[19152] = 8'hcb ;
            rom[19153] = 8'hf9 ;
            rom[19154] = 8'he5 ;
            rom[19155] = 8'hf3 ;
            rom[19156] = 8'he5 ;
            rom[19157] = 8'h08 ;
            rom[19158] = 8'he1 ;
            rom[19159] = 8'hff ;
            rom[19160] = 8'hd9 ;
            rom[19161] = 8'h05 ;
            rom[19162] = 8'hfb ;
            rom[19163] = 8'h23 ;
            rom[19164] = 8'h0a ;
            rom[19165] = 8'h26 ;
            rom[19166] = 8'he6 ;
            rom[19167] = 8'hde ;
            rom[19168] = 8'hf8 ;
            rom[19169] = 8'h0b ;
            rom[19170] = 8'hca ;
            rom[19171] = 8'haf ;
            rom[19172] = 8'h1d ;
            rom[19173] = 8'h27 ;
            rom[19174] = 8'h1b ;
            rom[19175] = 8'hce ;
            rom[19176] = 8'h04 ;
            rom[19177] = 8'h0e ;
            rom[19178] = 8'h1d ;
            rom[19179] = 8'h26 ;
            rom[19180] = 8'hcc ;
            rom[19181] = 8'hf3 ;
            rom[19182] = 8'hdb ;
            rom[19183] = 8'hfb ;
            rom[19184] = 8'h01 ;
            rom[19185] = 8'h2a ;
            rom[19186] = 8'h0f ;
            rom[19187] = 8'h3d ;
            rom[19188] = 8'h03 ;
            rom[19189] = 8'hf0 ;
            rom[19190] = 8'hf5 ;
            rom[19191] = 8'he0 ;
            rom[19192] = 8'hfc ;
            rom[19193] = 8'he1 ;
            rom[19194] = 8'h12 ;
            rom[19195] = 8'h1b ;
            rom[19196] = 8'h11 ;
            rom[19197] = 8'h13 ;
            rom[19198] = 8'h2a ;
            rom[19199] = 8'h07 ;
            rom[19200] = 8'he7 ;
            rom[19201] = 8'hf0 ;
            rom[19202] = 8'hd5 ;
            rom[19203] = 8'hf6 ;
            rom[19204] = 8'h11 ;
            rom[19205] = 8'hea ;
            rom[19206] = 8'h25 ;
            rom[19207] = 8'hd3 ;
            rom[19208] = 8'h0c ;
            rom[19209] = 8'hef ;
            rom[19210] = 8'he0 ;
            rom[19211] = 8'h00 ;
            rom[19212] = 8'h06 ;
            rom[19213] = 8'h0f ;
            rom[19214] = 8'haf ;
            rom[19215] = 8'h06 ;
            rom[19216] = 8'hee ;
            rom[19217] = 8'hf9 ;
            rom[19218] = 8'h24 ;
            rom[19219] = 8'hdc ;
            rom[19220] = 8'hd9 ;
            rom[19221] = 8'h14 ;
            rom[19222] = 8'h15 ;
            rom[19223] = 8'he8 ;
            rom[19224] = 8'he1 ;
            rom[19225] = 8'h04 ;
            rom[19226] = 8'hfe ;
            rom[19227] = 8'h04 ;
            rom[19228] = 8'hd3 ;
            rom[19229] = 8'hdb ;
            rom[19230] = 8'h0e ;
            rom[19231] = 8'h01 ;
            rom[19232] = 8'hf6 ;
            rom[19233] = 8'h02 ;
            rom[19234] = 8'hda ;
            rom[19235] = 8'h14 ;
            rom[19236] = 8'hd5 ;
            rom[19237] = 8'hf9 ;
            rom[19238] = 8'h21 ;
            rom[19239] = 8'he4 ;
            rom[19240] = 8'hf8 ;
            rom[19241] = 8'hf3 ;
            rom[19242] = 8'hfa ;
            rom[19243] = 8'h0a ;
            rom[19244] = 8'hdb ;
            rom[19245] = 8'h07 ;
            rom[19246] = 8'he8 ;
            rom[19247] = 8'h06 ;
            rom[19248] = 8'h14 ;
            rom[19249] = 8'hcf ;
            rom[19250] = 8'h0d ;
            rom[19251] = 8'h08 ;
            rom[19252] = 8'h01 ;
            rom[19253] = 8'hf8 ;
            rom[19254] = 8'hcf ;
            rom[19255] = 8'hfb ;
            rom[19256] = 8'hf0 ;
            rom[19257] = 8'h08 ;
            rom[19258] = 8'hf5 ;
            rom[19259] = 8'hec ;
            rom[19260] = 8'hf0 ;
            rom[19261] = 8'hea ;
            rom[19262] = 8'hf4 ;
            rom[19263] = 8'hf2 ;
            rom[19264] = 8'h17 ;
            rom[19265] = 8'hf9 ;
            rom[19266] = 8'hf5 ;
            rom[19267] = 8'h04 ;
            rom[19268] = 8'hfb ;
            rom[19269] = 8'hf5 ;
            rom[19270] = 8'heb ;
            rom[19271] = 8'hf4 ;
            rom[19272] = 8'hf2 ;
            rom[19273] = 8'hf1 ;
            rom[19274] = 8'h23 ;
            rom[19275] = 8'he9 ;
            rom[19276] = 8'h04 ;
            rom[19277] = 8'hdb ;
            rom[19278] = 8'hea ;
            rom[19279] = 8'h18 ;
            rom[19280] = 8'h11 ;
            rom[19281] = 8'h0a ;
            rom[19282] = 8'h01 ;
            rom[19283] = 8'h0a ;
            rom[19284] = 8'hf2 ;
            rom[19285] = 8'hd6 ;
            rom[19286] = 8'hf3 ;
            rom[19287] = 8'h12 ;
            rom[19288] = 8'hf4 ;
            rom[19289] = 8'h05 ;
            rom[19290] = 8'h17 ;
            rom[19291] = 8'h0d ;
            rom[19292] = 8'he7 ;
            rom[19293] = 8'h15 ;
            rom[19294] = 8'hf2 ;
            rom[19295] = 8'h05 ;
            rom[19296] = 8'hf7 ;
            rom[19297] = 8'he8 ;
            rom[19298] = 8'hbc ;
            rom[19299] = 8'hdf ;
            rom[19300] = 8'h0d ;
            rom[19301] = 8'h09 ;
            rom[19302] = 8'he8 ;
            rom[19303] = 8'hf4 ;
            rom[19304] = 8'hd8 ;
            rom[19305] = 8'hc2 ;
            rom[19306] = 8'hf6 ;
            rom[19307] = 8'h27 ;
            rom[19308] = 8'hf1 ;
            rom[19309] = 8'hee ;
            rom[19310] = 8'h09 ;
            rom[19311] = 8'h07 ;
            rom[19312] = 8'he3 ;
            rom[19313] = 8'h01 ;
            rom[19314] = 8'h0c ;
            rom[19315] = 8'h08 ;
            rom[19316] = 8'h0e ;
            rom[19317] = 8'h03 ;
            rom[19318] = 8'hd2 ;
            rom[19319] = 8'he4 ;
            rom[19320] = 8'h16 ;
            rom[19321] = 8'hf4 ;
            rom[19322] = 8'hd6 ;
            rom[19323] = 8'h24 ;
            rom[19324] = 8'h19 ;
            rom[19325] = 8'hf9 ;
            rom[19326] = 8'h14 ;
            rom[19327] = 8'h00 ;
            rom[19328] = 8'hf8 ;
            rom[19329] = 8'hfb ;
            rom[19330] = 8'h09 ;
            rom[19331] = 8'hf3 ;
            rom[19332] = 8'hcc ;
            rom[19333] = 8'hf4 ;
            rom[19334] = 8'h1d ;
            rom[19335] = 8'h28 ;
            rom[19336] = 8'h07 ;
            rom[19337] = 8'hff ;
            rom[19338] = 8'hfa ;
            rom[19339] = 8'hf3 ;
            rom[19340] = 8'h02 ;
            rom[19341] = 8'hea ;
            rom[19342] = 8'h13 ;
            rom[19343] = 8'h15 ;
            rom[19344] = 8'he3 ;
            rom[19345] = 8'he8 ;
            rom[19346] = 8'h0f ;
            rom[19347] = 8'he4 ;
            rom[19348] = 8'hf4 ;
            rom[19349] = 8'he4 ;
            rom[19350] = 8'heb ;
            rom[19351] = 8'h2c ;
            rom[19352] = 8'h07 ;
            rom[19353] = 8'h1e ;
            rom[19354] = 8'h09 ;
            rom[19355] = 8'hf4 ;
            rom[19356] = 8'he2 ;
            rom[19357] = 8'h15 ;
            rom[19358] = 8'h12 ;
            rom[19359] = 8'hf6 ;
            rom[19360] = 8'h0e ;
            rom[19361] = 8'hec ;
            rom[19362] = 8'h39 ;
            rom[19363] = 8'he3 ;
            rom[19364] = 8'hf3 ;
            rom[19365] = 8'hfb ;
            rom[19366] = 8'h22 ;
            rom[19367] = 8'hd3 ;
            rom[19368] = 8'h00 ;
            rom[19369] = 8'he8 ;
            rom[19370] = 8'h28 ;
            rom[19371] = 8'h09 ;
            rom[19372] = 8'h18 ;
            rom[19373] = 8'h08 ;
            rom[19374] = 8'hb6 ;
            rom[19375] = 8'h18 ;
            rom[19376] = 8'hef ;
            rom[19377] = 8'h18 ;
            rom[19378] = 8'h07 ;
            rom[19379] = 8'hd1 ;
            rom[19380] = 8'hfc ;
            rom[19381] = 8'hf8 ;
            rom[19382] = 8'hf2 ;
            rom[19383] = 8'h2f ;
            rom[19384] = 8'hf5 ;
            rom[19385] = 8'h07 ;
            rom[19386] = 8'hf0 ;
            rom[19387] = 8'hdf ;
            rom[19388] = 8'h1c ;
            rom[19389] = 8'h08 ;
            rom[19390] = 8'h18 ;
            rom[19391] = 8'h06 ;
            rom[19392] = 8'h12 ;
            rom[19393] = 8'h16 ;
            rom[19394] = 8'hf4 ;
            rom[19395] = 8'hf8 ;
            rom[19396] = 8'hfd ;
            rom[19397] = 8'h30 ;
            rom[19398] = 8'h0b ;
            rom[19399] = 8'h17 ;
            rom[19400] = 8'hc8 ;
            rom[19401] = 8'h2e ;
            rom[19402] = 8'hc5 ;
            rom[19403] = 8'hdb ;
            rom[19404] = 8'h1a ;
            rom[19405] = 8'h11 ;
            rom[19406] = 8'hf5 ;
            rom[19407] = 8'h0c ;
            rom[19408] = 8'h00 ;
            rom[19409] = 8'hf6 ;
            rom[19410] = 8'he8 ;
            rom[19411] = 8'h13 ;
            rom[19412] = 8'heb ;
            rom[19413] = 8'hdd ;
            rom[19414] = 8'hfe ;
            rom[19415] = 8'hf5 ;
            rom[19416] = 8'he7 ;
            rom[19417] = 8'h20 ;
            rom[19418] = 8'h18 ;
            rom[19419] = 8'hdc ;
            rom[19420] = 8'hf8 ;
            rom[19421] = 8'h0f ;
            rom[19422] = 8'h0f ;
            rom[19423] = 8'hf9 ;
            rom[19424] = 8'hef ;
            rom[19425] = 8'h29 ;
            rom[19426] = 8'hc5 ;
            rom[19427] = 8'h1f ;
            rom[19428] = 8'h17 ;
            rom[19429] = 8'h16 ;
            rom[19430] = 8'hfa ;
            rom[19431] = 8'h1a ;
            rom[19432] = 8'h10 ;
            rom[19433] = 8'hf4 ;
            rom[19434] = 8'hf4 ;
            rom[19435] = 8'h0e ;
            rom[19436] = 8'h06 ;
            rom[19437] = 8'hf1 ;
            rom[19438] = 8'hfe ;
            rom[19439] = 8'hfb ;
            rom[19440] = 8'hfa ;
            rom[19441] = 8'hcf ;
            rom[19442] = 8'h06 ;
            rom[19443] = 8'hfc ;
            rom[19444] = 8'h1d ;
            rom[19445] = 8'h20 ;
            rom[19446] = 8'h16 ;
            rom[19447] = 8'hdd ;
            rom[19448] = 8'hf5 ;
            rom[19449] = 8'h03 ;
            rom[19450] = 8'h0e ;
            rom[19451] = 8'hf1 ;
            rom[19452] = 8'h14 ;
            rom[19453] = 8'h01 ;
            rom[19454] = 8'h08 ;
            rom[19455] = 8'hf9 ;
            rom[19456] = 8'he7 ;
            rom[19457] = 8'hf4 ;
            rom[19458] = 8'hec ;
            rom[19459] = 8'hd4 ;
            rom[19460] = 8'h18 ;
            rom[19461] = 8'hfb ;
            rom[19462] = 8'hf9 ;
            rom[19463] = 8'h1a ;
            rom[19464] = 8'h13 ;
            rom[19465] = 8'heb ;
            rom[19466] = 8'h35 ;
            rom[19467] = 8'h10 ;
            rom[19468] = 8'h16 ;
            rom[19469] = 8'hf9 ;
            rom[19470] = 8'h01 ;
            rom[19471] = 8'h1a ;
            rom[19472] = 8'hcd ;
            rom[19473] = 8'h1d ;
            rom[19474] = 8'h0c ;
            rom[19475] = 8'h04 ;
            rom[19476] = 8'h0c ;
            rom[19477] = 8'h00 ;
            rom[19478] = 8'hd8 ;
            rom[19479] = 8'h25 ;
            rom[19480] = 8'hfb ;
            rom[19481] = 8'h0a ;
            rom[19482] = 8'h00 ;
            rom[19483] = 8'he4 ;
            rom[19484] = 8'h05 ;
            rom[19485] = 8'h31 ;
            rom[19486] = 8'h05 ;
            rom[19487] = 8'hed ;
            rom[19488] = 8'h0c ;
            rom[19489] = 8'hf1 ;
            rom[19490] = 8'h18 ;
            rom[19491] = 8'hff ;
            rom[19492] = 8'h1e ;
            rom[19493] = 8'h21 ;
            rom[19494] = 8'h1b ;
            rom[19495] = 8'he8 ;
            rom[19496] = 8'h16 ;
            rom[19497] = 8'h0b ;
            rom[19498] = 8'he6 ;
            rom[19499] = 8'h00 ;
            rom[19500] = 8'h09 ;
            rom[19501] = 8'h06 ;
            rom[19502] = 8'he3 ;
            rom[19503] = 8'he2 ;
            rom[19504] = 8'hf2 ;
            rom[19505] = 8'hf1 ;
            rom[19506] = 8'h0b ;
            rom[19507] = 8'h06 ;
            rom[19508] = 8'heb ;
            rom[19509] = 8'h0e ;
            rom[19510] = 8'h04 ;
            rom[19511] = 8'h02 ;
            rom[19512] = 8'hd4 ;
            rom[19513] = 8'hd8 ;
            rom[19514] = 8'h0c ;
            rom[19515] = 8'h04 ;
            rom[19516] = 8'h21 ;
            rom[19517] = 8'h0b ;
            rom[19518] = 8'h05 ;
            rom[19519] = 8'hfd ;
            rom[19520] = 8'hdb ;
            rom[19521] = 8'h11 ;
            rom[19522] = 8'h1c ;
            rom[19523] = 8'h0d ;
            rom[19524] = 8'hcd ;
            rom[19525] = 8'hfd ;
            rom[19526] = 8'h07 ;
            rom[19527] = 8'h02 ;
            rom[19528] = 8'he5 ;
            rom[19529] = 8'h0d ;
            rom[19530] = 8'hf0 ;
            rom[19531] = 8'h01 ;
            rom[19532] = 8'hef ;
            rom[19533] = 8'h02 ;
            rom[19534] = 8'h0a ;
            rom[19535] = 8'he5 ;
            rom[19536] = 8'h20 ;
            rom[19537] = 8'hfe ;
            rom[19538] = 8'hec ;
            rom[19539] = 8'hf1 ;
            rom[19540] = 8'hf2 ;
            rom[19541] = 8'h0b ;
            rom[19542] = 8'hf6 ;
            rom[19543] = 8'hf9 ;
            rom[19544] = 8'hf3 ;
            rom[19545] = 8'h02 ;
            rom[19546] = 8'hdc ;
            rom[19547] = 8'h05 ;
            rom[19548] = 8'hf0 ;
            rom[19549] = 8'hf6 ;
            rom[19550] = 8'h07 ;
            rom[19551] = 8'hff ;
            rom[19552] = 8'hec ;
            rom[19553] = 8'h13 ;
            rom[19554] = 8'hec ;
            rom[19555] = 8'hfc ;
            rom[19556] = 8'hf9 ;
            rom[19557] = 8'h09 ;
            rom[19558] = 8'h22 ;
            rom[19559] = 8'h16 ;
            rom[19560] = 8'hfd ;
            rom[19561] = 8'hf5 ;
            rom[19562] = 8'h39 ;
            rom[19563] = 8'h19 ;
            rom[19564] = 8'h06 ;
            rom[19565] = 8'hcb ;
            rom[19566] = 8'h10 ;
            rom[19567] = 8'hf3 ;
            rom[19568] = 8'hef ;
            rom[19569] = 8'hfd ;
            rom[19570] = 8'h35 ;
            rom[19571] = 8'h30 ;
            rom[19572] = 8'h46 ;
            rom[19573] = 8'h12 ;
            rom[19574] = 8'h09 ;
            rom[19575] = 8'h09 ;
            rom[19576] = 8'hff ;
            rom[19577] = 8'hf1 ;
            rom[19578] = 8'h16 ;
            rom[19579] = 8'hf0 ;
            rom[19580] = 8'h03 ;
            rom[19581] = 8'h12 ;
            rom[19582] = 8'h0f ;
            rom[19583] = 8'he2 ;
            rom[19584] = 8'hd4 ;
            rom[19585] = 8'hfc ;
            rom[19586] = 8'h25 ;
            rom[19587] = 8'h07 ;
            rom[19588] = 8'hec ;
            rom[19589] = 8'h23 ;
            rom[19590] = 8'h05 ;
            rom[19591] = 8'hff ;
            rom[19592] = 8'h20 ;
            rom[19593] = 8'hf1 ;
            rom[19594] = 8'h2a ;
            rom[19595] = 8'hdd ;
            rom[19596] = 8'h11 ;
            rom[19597] = 8'h08 ;
            rom[19598] = 8'hfb ;
            rom[19599] = 8'hfb ;
            rom[19600] = 8'hdb ;
            rom[19601] = 8'hde ;
            rom[19602] = 8'h1a ;
            rom[19603] = 8'he9 ;
            rom[19604] = 8'hea ;
            rom[19605] = 8'h09 ;
            rom[19606] = 8'h04 ;
            rom[19607] = 8'h05 ;
            rom[19608] = 8'hf1 ;
            rom[19609] = 8'h14 ;
            rom[19610] = 8'hf4 ;
            rom[19611] = 8'he4 ;
            rom[19612] = 8'h07 ;
            rom[19613] = 8'he9 ;
            rom[19614] = 8'h0b ;
            rom[19615] = 8'hd2 ;
            rom[19616] = 8'hd6 ;
            rom[19617] = 8'hcc ;
            rom[19618] = 8'h0b ;
            rom[19619] = 8'h15 ;
            rom[19620] = 8'hc2 ;
            rom[19621] = 8'h0c ;
            rom[19622] = 8'h12 ;
            rom[19623] = 8'h10 ;
            rom[19624] = 8'he9 ;
            rom[19625] = 8'hfc ;
            rom[19626] = 8'h18 ;
            rom[19627] = 8'h1e ;
            rom[19628] = 8'h05 ;
            rom[19629] = 8'he3 ;
            rom[19630] = 8'h29 ;
            rom[19631] = 8'he9 ;
            rom[19632] = 8'h2b ;
            rom[19633] = 8'he4 ;
            rom[19634] = 8'h01 ;
            rom[19635] = 8'h18 ;
            rom[19636] = 8'he2 ;
            rom[19637] = 8'hea ;
            rom[19638] = 8'h1f ;
            rom[19639] = 8'h3a ;
            rom[19640] = 8'h08 ;
            rom[19641] = 8'hf0 ;
            rom[19642] = 8'h13 ;
            rom[19643] = 8'h05 ;
            rom[19644] = 8'h34 ;
            rom[19645] = 8'hf9 ;
            rom[19646] = 8'hf5 ;
            rom[19647] = 8'h34 ;
            rom[19648] = 8'h0b ;
            rom[19649] = 8'hd5 ;
            rom[19650] = 8'he4 ;
            rom[19651] = 8'h0d ;
            rom[19652] = 8'he8 ;
            rom[19653] = 8'h14 ;
            rom[19654] = 8'h0d ;
            rom[19655] = 8'he1 ;
            rom[19656] = 8'h01 ;
            rom[19657] = 8'h15 ;
            rom[19658] = 8'hf5 ;
            rom[19659] = 8'hea ;
            rom[19660] = 8'hf5 ;
            rom[19661] = 8'h03 ;
            rom[19662] = 8'he2 ;
            rom[19663] = 8'h21 ;
            rom[19664] = 8'hff ;
            rom[19665] = 8'hf2 ;
            rom[19666] = 8'hf4 ;
            rom[19667] = 8'hff ;
            rom[19668] = 8'hf2 ;
            rom[19669] = 8'h0e ;
            rom[19670] = 8'hd7 ;
            rom[19671] = 8'h1e ;
            rom[19672] = 8'hf2 ;
            rom[19673] = 8'he7 ;
            rom[19674] = 8'hdb ;
            rom[19675] = 8'he0 ;
            rom[19676] = 8'h01 ;
            rom[19677] = 8'h1b ;
            rom[19678] = 8'he6 ;
            rom[19679] = 8'h24 ;
            rom[19680] = 8'hf2 ;
            rom[19681] = 8'h05 ;
            rom[19682] = 8'h09 ;
            rom[19683] = 8'hfd ;
            rom[19684] = 8'hf8 ;
            rom[19685] = 8'h14 ;
            rom[19686] = 8'h13 ;
            rom[19687] = 8'h09 ;
            rom[19688] = 8'hea ;
            rom[19689] = 8'hf8 ;
            rom[19690] = 8'hdf ;
            rom[19691] = 8'hdf ;
            rom[19692] = 8'h0f ;
            rom[19693] = 8'he6 ;
            rom[19694] = 8'h17 ;
            rom[19695] = 8'h03 ;
            rom[19696] = 8'h1b ;
            rom[19697] = 8'hf1 ;
            rom[19698] = 8'h0f ;
            rom[19699] = 8'h0c ;
            rom[19700] = 8'h2a ;
            rom[19701] = 8'h07 ;
            rom[19702] = 8'hea ;
            rom[19703] = 8'hf5 ;
            rom[19704] = 8'hf7 ;
            rom[19705] = 8'h03 ;
            rom[19706] = 8'hef ;
            rom[19707] = 8'h16 ;
            rom[19708] = 8'h07 ;
            rom[19709] = 8'hd1 ;
            rom[19710] = 8'h2a ;
            rom[19711] = 8'hf1 ;
            rom[19712] = 8'hf4 ;
            rom[19713] = 8'h03 ;
            rom[19714] = 8'h0f ;
            rom[19715] = 8'hdb ;
            rom[19716] = 8'h0b ;
            rom[19717] = 8'hfe ;
            rom[19718] = 8'hde ;
            rom[19719] = 8'h11 ;
            rom[19720] = 8'h29 ;
            rom[19721] = 8'h0f ;
            rom[19722] = 8'hdd ;
            rom[19723] = 8'h0d ;
            rom[19724] = 8'he8 ;
            rom[19725] = 8'hed ;
            rom[19726] = 8'h21 ;
            rom[19727] = 8'h14 ;
            rom[19728] = 8'hf7 ;
            rom[19729] = 8'hf8 ;
            rom[19730] = 8'h06 ;
            rom[19731] = 8'h10 ;
            rom[19732] = 8'h19 ;
            rom[19733] = 8'hd8 ;
            rom[19734] = 8'hf6 ;
            rom[19735] = 8'h10 ;
            rom[19736] = 8'h25 ;
            rom[19737] = 8'hf2 ;
            rom[19738] = 8'hfb ;
            rom[19739] = 8'hf2 ;
            rom[19740] = 8'h15 ;
            rom[19741] = 8'h2c ;
            rom[19742] = 8'h1c ;
            rom[19743] = 8'he2 ;
            rom[19744] = 8'hf5 ;
            rom[19745] = 8'hee ;
            rom[19746] = 8'h17 ;
            rom[19747] = 8'hf6 ;
            rom[19748] = 8'h0b ;
            rom[19749] = 8'h05 ;
            rom[19750] = 8'h2b ;
            rom[19751] = 8'hea ;
            rom[19752] = 8'he3 ;
            rom[19753] = 8'he5 ;
            rom[19754] = 8'h05 ;
            rom[19755] = 8'hfe ;
            rom[19756] = 8'hfc ;
            rom[19757] = 8'h0a ;
            rom[19758] = 8'hf5 ;
            rom[19759] = 8'hf2 ;
            rom[19760] = 8'h0b ;
            rom[19761] = 8'he5 ;
            rom[19762] = 8'h0e ;
            rom[19763] = 8'hf1 ;
            rom[19764] = 8'hf5 ;
            rom[19765] = 8'hf6 ;
            rom[19766] = 8'h15 ;
            rom[19767] = 8'hf8 ;
            rom[19768] = 8'h10 ;
            rom[19769] = 8'h01 ;
            rom[19770] = 8'he0 ;
            rom[19771] = 8'hd9 ;
            rom[19772] = 8'hff ;
            rom[19773] = 8'hec ;
            rom[19774] = 8'h0d ;
            rom[19775] = 8'hef ;
            rom[19776] = 8'hf4 ;
            rom[19777] = 8'h33 ;
            rom[19778] = 8'h30 ;
            rom[19779] = 8'h2a ;
            rom[19780] = 8'hf4 ;
            rom[19781] = 8'hf4 ;
            rom[19782] = 8'h2a ;
            rom[19783] = 8'h00 ;
            rom[19784] = 8'hd1 ;
            rom[19785] = 8'h1e ;
            rom[19786] = 8'he9 ;
            rom[19787] = 8'he3 ;
            rom[19788] = 8'hef ;
            rom[19789] = 8'h0e ;
            rom[19790] = 8'h09 ;
            rom[19791] = 8'hef ;
            rom[19792] = 8'h0f ;
            rom[19793] = 8'h14 ;
            rom[19794] = 8'hec ;
            rom[19795] = 8'hfa ;
            rom[19796] = 8'hec ;
            rom[19797] = 8'h0d ;
            rom[19798] = 8'h0b ;
            rom[19799] = 8'he1 ;
            rom[19800] = 8'hfa ;
            rom[19801] = 8'h06 ;
            rom[19802] = 8'h08 ;
            rom[19803] = 8'hfe ;
            rom[19804] = 8'hfb ;
            rom[19805] = 8'hf7 ;
            rom[19806] = 8'h06 ;
            rom[19807] = 8'hee ;
            rom[19808] = 8'h02 ;
            rom[19809] = 8'h09 ;
            rom[19810] = 8'hf2 ;
            rom[19811] = 8'hed ;
            rom[19812] = 8'hfe ;
            rom[19813] = 8'h01 ;
            rom[19814] = 8'he4 ;
            rom[19815] = 8'hfe ;
            rom[19816] = 8'h12 ;
            rom[19817] = 8'hfa ;
            rom[19818] = 8'h36 ;
            rom[19819] = 8'hf0 ;
            rom[19820] = 8'h04 ;
            rom[19821] = 8'he9 ;
            rom[19822] = 8'h01 ;
            rom[19823] = 8'hf4 ;
            rom[19824] = 8'hf8 ;
            rom[19825] = 8'hdc ;
            rom[19826] = 8'hea ;
            rom[19827] = 8'h27 ;
            rom[19828] = 8'h09 ;
            rom[19829] = 8'h1e ;
            rom[19830] = 8'hfd ;
            rom[19831] = 8'hc9 ;
            rom[19832] = 8'hf6 ;
            rom[19833] = 8'hf8 ;
            rom[19834] = 8'h13 ;
            rom[19835] = 8'h1b ;
            rom[19836] = 8'hed ;
            rom[19837] = 8'hff ;
            rom[19838] = 8'hfb ;
            rom[19839] = 8'h1b ;
            rom[19840] = 8'hcd ;
            rom[19841] = 8'hfb ;
            rom[19842] = 8'h06 ;
            rom[19843] = 8'he1 ;
            rom[19844] = 8'h1b ;
            rom[19845] = 8'hf5 ;
            rom[19846] = 8'heb ;
            rom[19847] = 8'hdf ;
            rom[19848] = 8'hfa ;
            rom[19849] = 8'he1 ;
            rom[19850] = 8'h0a ;
            rom[19851] = 8'he3 ;
            rom[19852] = 8'hf1 ;
            rom[19853] = 8'h35 ;
            rom[19854] = 8'hd5 ;
            rom[19855] = 8'h13 ;
            rom[19856] = 8'h1e ;
            rom[19857] = 8'h05 ;
            rom[19858] = 8'hf0 ;
            rom[19859] = 8'hc8 ;
            rom[19860] = 8'he4 ;
            rom[19861] = 8'hfb ;
            rom[19862] = 8'h45 ;
            rom[19863] = 8'hec ;
            rom[19864] = 8'h2f ;
            rom[19865] = 8'h23 ;
            rom[19866] = 8'hc8 ;
            rom[19867] = 8'h2b ;
            rom[19868] = 8'hf1 ;
            rom[19869] = 8'h11 ;
            rom[19870] = 8'h21 ;
            rom[19871] = 8'h1b ;
            rom[19872] = 8'h13 ;
            rom[19873] = 8'hff ;
            rom[19874] = 8'hdf ;
            rom[19875] = 8'hf2 ;
            rom[19876] = 8'he0 ;
            rom[19877] = 8'hc7 ;
            rom[19878] = 8'h18 ;
            rom[19879] = 8'hf7 ;
            rom[19880] = 8'he6 ;
            rom[19881] = 8'hd2 ;
            rom[19882] = 8'hef ;
            rom[19883] = 8'h10 ;
            rom[19884] = 8'h04 ;
            rom[19885] = 8'he2 ;
            rom[19886] = 8'h13 ;
            rom[19887] = 8'hf9 ;
            rom[19888] = 8'h0d ;
            rom[19889] = 8'h04 ;
            rom[19890] = 8'hee ;
            rom[19891] = 8'hf6 ;
            rom[19892] = 8'he6 ;
            rom[19893] = 8'hef ;
            rom[19894] = 8'h14 ;
            rom[19895] = 8'h04 ;
            rom[19896] = 8'h08 ;
            rom[19897] = 8'hf4 ;
            rom[19898] = 8'heb ;
            rom[19899] = 8'hef ;
            rom[19900] = 8'h08 ;
            rom[19901] = 8'he8 ;
            rom[19902] = 8'hfc ;
            rom[19903] = 8'h02 ;
            rom[19904] = 8'h0a ;
            rom[19905] = 8'hfd ;
            rom[19906] = 8'hfe ;
            rom[19907] = 8'h1a ;
            rom[19908] = 8'h0b ;
            rom[19909] = 8'he3 ;
            rom[19910] = 8'hf1 ;
            rom[19911] = 8'he9 ;
            rom[19912] = 8'h06 ;
            rom[19913] = 8'hee ;
            rom[19914] = 8'hd3 ;
            rom[19915] = 8'hed ;
            rom[19916] = 8'hd9 ;
            rom[19917] = 8'hb1 ;
            rom[19918] = 8'hdb ;
            rom[19919] = 8'h1a ;
            rom[19920] = 8'h00 ;
            rom[19921] = 8'h3f ;
            rom[19922] = 8'h05 ;
            rom[19923] = 8'he6 ;
            rom[19924] = 8'h18 ;
            rom[19925] = 8'h11 ;
            rom[19926] = 8'hcd ;
            rom[19927] = 8'h25 ;
            rom[19928] = 8'hea ;
            rom[19929] = 8'hed ;
            rom[19930] = 8'hd8 ;
            rom[19931] = 8'hf9 ;
            rom[19932] = 8'hfe ;
            rom[19933] = 8'h0c ;
            rom[19934] = 8'hbe ;
            rom[19935] = 8'hdb ;
            rom[19936] = 8'hf6 ;
            rom[19937] = 8'h2a ;
            rom[19938] = 8'h03 ;
            rom[19939] = 8'hf0 ;
            rom[19940] = 8'h04 ;
            rom[19941] = 8'hf5 ;
            rom[19942] = 8'h0c ;
            rom[19943] = 8'hd8 ;
            rom[19944] = 8'h0b ;
            rom[19945] = 8'h02 ;
            rom[19946] = 8'he0 ;
            rom[19947] = 8'h12 ;
            rom[19948] = 8'h04 ;
            rom[19949] = 8'hfd ;
            rom[19950] = 8'hf3 ;
            rom[19951] = 8'h23 ;
            rom[19952] = 8'hfb ;
            rom[19953] = 8'h06 ;
            rom[19954] = 8'h1b ;
            rom[19955] = 8'h0c ;
            rom[19956] = 8'heb ;
            rom[19957] = 8'he8 ;
            rom[19958] = 8'h04 ;
            rom[19959] = 8'h07 ;
            rom[19960] = 8'hf9 ;
            rom[19961] = 8'hfb ;
            rom[19962] = 8'had ;
            rom[19963] = 8'hf2 ;
            rom[19964] = 8'h0a ;
            rom[19965] = 8'h0d ;
            rom[19966] = 8'h07 ;
            rom[19967] = 8'h0d ;
            rom[19968] = 8'h04 ;
            rom[19969] = 8'hec ;
            rom[19970] = 8'h0f ;
            rom[19971] = 8'h03 ;
            rom[19972] = 8'hf4 ;
            rom[19973] = 8'h28 ;
            rom[19974] = 8'hff ;
            rom[19975] = 8'h0b ;
            rom[19976] = 8'hf9 ;
            rom[19977] = 8'hfe ;
            rom[19978] = 8'h0e ;
            rom[19979] = 8'hfd ;
            rom[19980] = 8'he0 ;
            rom[19981] = 8'h10 ;
            rom[19982] = 8'h2e ;
            rom[19983] = 8'he0 ;
            rom[19984] = 8'h12 ;
            rom[19985] = 8'h0c ;
            rom[19986] = 8'hf8 ;
            rom[19987] = 8'h06 ;
            rom[19988] = 8'h05 ;
            rom[19989] = 8'hd0 ;
            rom[19990] = 8'h06 ;
            rom[19991] = 8'h13 ;
            rom[19992] = 8'hf1 ;
            rom[19993] = 8'h0a ;
            rom[19994] = 8'he5 ;
            rom[19995] = 8'hba ;
            rom[19996] = 8'hc8 ;
            rom[19997] = 8'h10 ;
            rom[19998] = 8'h0f ;
            rom[19999] = 8'h0b ;
            rom[20000] = 8'h18 ;
            rom[20001] = 8'hdd ;
            rom[20002] = 8'hf6 ;
            rom[20003] = 8'hf3 ;
            rom[20004] = 8'hf8 ;
            rom[20005] = 8'he4 ;
            rom[20006] = 8'h0d ;
            rom[20007] = 8'he7 ;
            rom[20008] = 8'hde ;
            rom[20009] = 8'hc4 ;
            rom[20010] = 8'hf4 ;
            rom[20011] = 8'h22 ;
            rom[20012] = 8'h09 ;
            rom[20013] = 8'hec ;
            rom[20014] = 8'hfc ;
            rom[20015] = 8'h05 ;
            rom[20016] = 8'hc3 ;
            rom[20017] = 8'he3 ;
            rom[20018] = 8'he9 ;
            rom[20019] = 8'h17 ;
            rom[20020] = 8'hf8 ;
            rom[20021] = 8'hd7 ;
            rom[20022] = 8'heb ;
            rom[20023] = 8'h03 ;
            rom[20024] = 8'hf3 ;
            rom[20025] = 8'heb ;
            rom[20026] = 8'h23 ;
            rom[20027] = 8'h13 ;
            rom[20028] = 8'hf3 ;
            rom[20029] = 8'hef ;
            rom[20030] = 8'hf6 ;
            rom[20031] = 8'h21 ;
            rom[20032] = 8'h02 ;
            rom[20033] = 8'h0f ;
            rom[20034] = 8'hec ;
            rom[20035] = 8'hd2 ;
            rom[20036] = 8'h09 ;
            rom[20037] = 8'hd3 ;
            rom[20038] = 8'h23 ;
            rom[20039] = 8'he7 ;
            rom[20040] = 8'h2c ;
            rom[20041] = 8'h00 ;
            rom[20042] = 8'hf1 ;
            rom[20043] = 8'h08 ;
            rom[20044] = 8'he4 ;
            rom[20045] = 8'hdf ;
            rom[20046] = 8'h0c ;
            rom[20047] = 8'h04 ;
            rom[20048] = 8'h00 ;
            rom[20049] = 8'h27 ;
            rom[20050] = 8'hfd ;
            rom[20051] = 8'hce ;
            rom[20052] = 8'he9 ;
            rom[20053] = 8'h2e ;
            rom[20054] = 8'h26 ;
            rom[20055] = 8'h0a ;
            rom[20056] = 8'h30 ;
            rom[20057] = 8'hd1 ;
            rom[20058] = 8'he5 ;
            rom[20059] = 8'h01 ;
            rom[20060] = 8'hee ;
            rom[20061] = 8'h0b ;
            rom[20062] = 8'hf4 ;
            rom[20063] = 8'hf4 ;
            rom[20064] = 8'hef ;
            rom[20065] = 8'hff ;
            rom[20066] = 8'h18 ;
            rom[20067] = 8'hf8 ;
            rom[20068] = 8'heb ;
            rom[20069] = 8'hd3 ;
            rom[20070] = 8'hf1 ;
            rom[20071] = 8'hfa ;
            rom[20072] = 8'hff ;
            rom[20073] = 8'hf0 ;
            rom[20074] = 8'hf0 ;
            rom[20075] = 8'h02 ;
            rom[20076] = 8'h28 ;
            rom[20077] = 8'he3 ;
            rom[20078] = 8'h12 ;
            rom[20079] = 8'hf9 ;
            rom[20080] = 8'hdb ;
            rom[20081] = 8'hd6 ;
            rom[20082] = 8'h11 ;
            rom[20083] = 8'h10 ;
            rom[20084] = 8'h08 ;
            rom[20085] = 8'h11 ;
            rom[20086] = 8'hed ;
            rom[20087] = 8'hfc ;
            rom[20088] = 8'hec ;
            rom[20089] = 8'hfe ;
            rom[20090] = 8'hf4 ;
            rom[20091] = 8'hee ;
            rom[20092] = 8'hcf ;
            rom[20093] = 8'h03 ;
            rom[20094] = 8'hed ;
            rom[20095] = 8'h0e ;
            rom[20096] = 8'hfb ;
            rom[20097] = 8'hf9 ;
            rom[20098] = 8'hd6 ;
            rom[20099] = 8'h11 ;
            rom[20100] = 8'h05 ;
            rom[20101] = 8'h11 ;
            rom[20102] = 8'hf3 ;
            rom[20103] = 8'h08 ;
            rom[20104] = 8'hfe ;
            rom[20105] = 8'hf4 ;
            rom[20106] = 8'h0b ;
            rom[20107] = 8'hfa ;
            rom[20108] = 8'hcb ;
            rom[20109] = 8'h0d ;
            rom[20110] = 8'h22 ;
            rom[20111] = 8'h26 ;
            rom[20112] = 8'h00 ;
            rom[20113] = 8'h03 ;
            rom[20114] = 8'hf7 ;
            rom[20115] = 8'he4 ;
            rom[20116] = 8'h19 ;
            rom[20117] = 8'hec ;
            rom[20118] = 8'hdd ;
            rom[20119] = 8'hce ;
            rom[20120] = 8'hd0 ;
            rom[20121] = 8'h20 ;
            rom[20122] = 8'h05 ;
            rom[20123] = 8'hdb ;
            rom[20124] = 8'h18 ;
            rom[20125] = 8'he1 ;
            rom[20126] = 8'h10 ;
            rom[20127] = 8'hee ;
            rom[20128] = 8'h01 ;
            rom[20129] = 8'hf8 ;
            rom[20130] = 8'hea ;
            rom[20131] = 8'hd8 ;
            rom[20132] = 8'hdc ;
            rom[20133] = 8'h15 ;
            rom[20134] = 8'hf7 ;
            rom[20135] = 8'he9 ;
            rom[20136] = 8'hcf ;
            rom[20137] = 8'h01 ;
            rom[20138] = 8'hfe ;
            rom[20139] = 8'h02 ;
            rom[20140] = 8'h1d ;
            rom[20141] = 8'hfa ;
            rom[20142] = 8'he4 ;
            rom[20143] = 8'h08 ;
            rom[20144] = 8'h0e ;
            rom[20145] = 8'hc6 ;
            rom[20146] = 8'hc6 ;
            rom[20147] = 8'h22 ;
            rom[20148] = 8'hd2 ;
            rom[20149] = 8'hff ;
            rom[20150] = 8'h15 ;
            rom[20151] = 8'h0e ;
            rom[20152] = 8'hfb ;
            rom[20153] = 8'he3 ;
            rom[20154] = 8'hf2 ;
            rom[20155] = 8'h22 ;
            rom[20156] = 8'h0f ;
            rom[20157] = 8'h05 ;
            rom[20158] = 8'hfb ;
            rom[20159] = 8'hf7 ;
            rom[20160] = 8'h29 ;
            rom[20161] = 8'he8 ;
            rom[20162] = 8'h05 ;
            rom[20163] = 8'he4 ;
            rom[20164] = 8'hff ;
            rom[20165] = 8'hf9 ;
            rom[20166] = 8'hfc ;
            rom[20167] = 8'hf8 ;
            rom[20168] = 8'hf6 ;
            rom[20169] = 8'hec ;
            rom[20170] = 8'h08 ;
            rom[20171] = 8'he5 ;
            rom[20172] = 8'hf4 ;
            rom[20173] = 8'hdf ;
            rom[20174] = 8'h0b ;
            rom[20175] = 8'hff ;
            rom[20176] = 8'h17 ;
            rom[20177] = 8'hf2 ;
            rom[20178] = 8'h03 ;
            rom[20179] = 8'hd7 ;
            rom[20180] = 8'hda ;
            rom[20181] = 8'h08 ;
            rom[20182] = 8'hf7 ;
            rom[20183] = 8'h10 ;
            rom[20184] = 8'h06 ;
            rom[20185] = 8'hf4 ;
            rom[20186] = 8'hf0 ;
            rom[20187] = 8'hef ;
            rom[20188] = 8'hb8 ;
            rom[20189] = 8'h22 ;
            rom[20190] = 8'hca ;
            rom[20191] = 8'h06 ;
            rom[20192] = 8'he5 ;
            rom[20193] = 8'hec ;
            rom[20194] = 8'he4 ;
            rom[20195] = 8'hd6 ;
            rom[20196] = 8'h19 ;
            rom[20197] = 8'hfa ;
            rom[20198] = 8'h0a ;
            rom[20199] = 8'hde ;
            rom[20200] = 8'h04 ;
            rom[20201] = 8'he0 ;
            rom[20202] = 8'he4 ;
            rom[20203] = 8'he0 ;
            rom[20204] = 8'h01 ;
            rom[20205] = 8'hdc ;
            rom[20206] = 8'hdf ;
            rom[20207] = 8'hfd ;
            rom[20208] = 8'h01 ;
            rom[20209] = 8'hf4 ;
            rom[20210] = 8'h16 ;
            rom[20211] = 8'hfb ;
            rom[20212] = 8'h14 ;
            rom[20213] = 8'h19 ;
            rom[20214] = 8'h07 ;
            rom[20215] = 8'hef ;
            rom[20216] = 8'hc6 ;
            rom[20217] = 8'he8 ;
            rom[20218] = 8'h09 ;
            rom[20219] = 8'he7 ;
            rom[20220] = 8'hff ;
            rom[20221] = 8'h13 ;
            rom[20222] = 8'hf1 ;
            rom[20223] = 8'h08 ;
            rom[20224] = 8'hfd ;
            rom[20225] = 8'he0 ;
            rom[20226] = 8'hf8 ;
            rom[20227] = 8'h0d ;
            rom[20228] = 8'h03 ;
            rom[20229] = 8'h07 ;
            rom[20230] = 8'h01 ;
            rom[20231] = 8'he7 ;
            rom[20232] = 8'h07 ;
            rom[20233] = 8'hd6 ;
            rom[20234] = 8'h1b ;
            rom[20235] = 8'heb ;
            rom[20236] = 8'hf0 ;
            rom[20237] = 8'h0a ;
            rom[20238] = 8'h00 ;
            rom[20239] = 8'h0e ;
            rom[20240] = 8'h0f ;
            rom[20241] = 8'h24 ;
            rom[20242] = 8'hef ;
            rom[20243] = 8'hda ;
            rom[20244] = 8'h28 ;
            rom[20245] = 8'h31 ;
            rom[20246] = 8'hed ;
            rom[20247] = 8'hf7 ;
            rom[20248] = 8'hf0 ;
            rom[20249] = 8'h23 ;
            rom[20250] = 8'h04 ;
            rom[20251] = 8'hf4 ;
            rom[20252] = 8'h0c ;
            rom[20253] = 8'h07 ;
            rom[20254] = 8'h21 ;
            rom[20255] = 8'h12 ;
            rom[20256] = 8'h14 ;
            rom[20257] = 8'h0b ;
            rom[20258] = 8'he4 ;
            rom[20259] = 8'hbf ;
            rom[20260] = 8'hfe ;
            rom[20261] = 8'hfe ;
            rom[20262] = 8'h0f ;
            rom[20263] = 8'h12 ;
            rom[20264] = 8'h00 ;
            rom[20265] = 8'h07 ;
            rom[20266] = 8'h07 ;
            rom[20267] = 8'hfd ;
            rom[20268] = 8'h0c ;
            rom[20269] = 8'hf9 ;
            rom[20270] = 8'hf5 ;
            rom[20271] = 8'hfe ;
            rom[20272] = 8'he3 ;
            rom[20273] = 8'he4 ;
            rom[20274] = 8'he1 ;
            rom[20275] = 8'h09 ;
            rom[20276] = 8'hd4 ;
            rom[20277] = 8'h00 ;
            rom[20278] = 8'h03 ;
            rom[20279] = 8'hd7 ;
            rom[20280] = 8'hef ;
            rom[20281] = 8'hf5 ;
            rom[20282] = 8'h0f ;
            rom[20283] = 8'hf7 ;
            rom[20284] = 8'h1c ;
            rom[20285] = 8'hf4 ;
            rom[20286] = 8'hf1 ;
            rom[20287] = 8'h01 ;
            rom[20288] = 8'hf7 ;
            rom[20289] = 8'hd2 ;
            rom[20290] = 8'hf8 ;
            rom[20291] = 8'h07 ;
            rom[20292] = 8'h1c ;
            rom[20293] = 8'hf3 ;
            rom[20294] = 8'hfc ;
            rom[20295] = 8'h0e ;
            rom[20296] = 8'h1e ;
            rom[20297] = 8'h0c ;
            rom[20298] = 8'h06 ;
            rom[20299] = 8'h1c ;
            rom[20300] = 8'h20 ;
            rom[20301] = 8'hd7 ;
            rom[20302] = 8'hdc ;
            rom[20303] = 8'h0f ;
            rom[20304] = 8'hda ;
            rom[20305] = 8'hf4 ;
            rom[20306] = 8'hfa ;
            rom[20307] = 8'hdc ;
            rom[20308] = 8'hec ;
            rom[20309] = 8'h00 ;
            rom[20310] = 8'hef ;
            rom[20311] = 8'h26 ;
            rom[20312] = 8'hed ;
            rom[20313] = 8'hea ;
            rom[20314] = 8'hf4 ;
            rom[20315] = 8'hf5 ;
            rom[20316] = 8'he8 ;
            rom[20317] = 8'h29 ;
            rom[20318] = 8'hfd ;
            rom[20319] = 8'h00 ;
            rom[20320] = 8'hf5 ;
            rom[20321] = 8'h04 ;
            rom[20322] = 8'hee ;
            rom[20323] = 8'hcd ;
            rom[20324] = 8'hf9 ;
            rom[20325] = 8'h02 ;
            rom[20326] = 8'h27 ;
            rom[20327] = 8'hd9 ;
            rom[20328] = 8'h00 ;
            rom[20329] = 8'h18 ;
            rom[20330] = 8'h01 ;
            rom[20331] = 8'h12 ;
            rom[20332] = 8'h0d ;
            rom[20333] = 8'hf1 ;
            rom[20334] = 8'he1 ;
            rom[20335] = 8'h10 ;
            rom[20336] = 8'h23 ;
            rom[20337] = 8'h23 ;
            rom[20338] = 8'h41 ;
            rom[20339] = 8'h0c ;
            rom[20340] = 8'hf6 ;
            rom[20341] = 8'he5 ;
            rom[20342] = 8'hfa ;
            rom[20343] = 8'h0c ;
            rom[20344] = 8'hd5 ;
            rom[20345] = 8'h22 ;
            rom[20346] = 8'h09 ;
            rom[20347] = 8'hf2 ;
            rom[20348] = 8'h06 ;
            rom[20349] = 8'hfe ;
            rom[20350] = 8'h13 ;
            rom[20351] = 8'h20 ;
            rom[20352] = 8'hf9 ;
            rom[20353] = 8'h02 ;
            rom[20354] = 8'h02 ;
            rom[20355] = 8'h00 ;
            rom[20356] = 8'h06 ;
            rom[20357] = 8'hfd ;
            rom[20358] = 8'hdc ;
            rom[20359] = 8'he0 ;
            rom[20360] = 8'hcd ;
            rom[20361] = 8'h10 ;
            rom[20362] = 8'he6 ;
            rom[20363] = 8'hed ;
            rom[20364] = 8'h02 ;
            rom[20365] = 8'hf8 ;
            rom[20366] = 8'hfa ;
            rom[20367] = 8'hd8 ;
            rom[20368] = 8'h22 ;
            rom[20369] = 8'hf9 ;
            rom[20370] = 8'hed ;
            rom[20371] = 8'h15 ;
            rom[20372] = 8'h0c ;
            rom[20373] = 8'h07 ;
            rom[20374] = 8'h04 ;
            rom[20375] = 8'hd4 ;
            rom[20376] = 8'hde ;
            rom[20377] = 8'h0c ;
            rom[20378] = 8'hf6 ;
            rom[20379] = 8'hdd ;
            rom[20380] = 8'hec ;
            rom[20381] = 8'hd3 ;
            rom[20382] = 8'he1 ;
            rom[20383] = 8'h12 ;
            rom[20384] = 8'hbe ;
            rom[20385] = 8'hea ;
            rom[20386] = 8'hde ;
            rom[20387] = 8'h01 ;
            rom[20388] = 8'h0f ;
            rom[20389] = 8'he3 ;
            rom[20390] = 8'hff ;
            rom[20391] = 8'heb ;
            rom[20392] = 8'hee ;
            rom[20393] = 8'hd7 ;
            rom[20394] = 8'hd3 ;
            rom[20395] = 8'hf4 ;
            rom[20396] = 8'he8 ;
            rom[20397] = 8'h08 ;
            rom[20398] = 8'hd4 ;
            rom[20399] = 8'he9 ;
            rom[20400] = 8'h10 ;
            rom[20401] = 8'hfe ;
            rom[20402] = 8'h00 ;
            rom[20403] = 8'h08 ;
            rom[20404] = 8'h04 ;
            rom[20405] = 8'hef ;
            rom[20406] = 8'hd1 ;
            rom[20407] = 8'hed ;
            rom[20408] = 8'h05 ;
            rom[20409] = 8'h02 ;
            rom[20410] = 8'hf0 ;
            rom[20411] = 8'hfd ;
            rom[20412] = 8'hd4 ;
            rom[20413] = 8'hd4 ;
            rom[20414] = 8'hf7 ;
            rom[20415] = 8'hea ;
            rom[20416] = 8'h36 ;
            rom[20417] = 8'hf2 ;
            rom[20418] = 8'h0e ;
            rom[20419] = 8'hf2 ;
            rom[20420] = 8'h0e ;
            rom[20421] = 8'hdb ;
            rom[20422] = 8'he5 ;
            rom[20423] = 8'hf2 ;
            rom[20424] = 8'h09 ;
            rom[20425] = 8'hed ;
            rom[20426] = 8'hf8 ;
            rom[20427] = 8'h00 ;
            rom[20428] = 8'he8 ;
            rom[20429] = 8'hef ;
            rom[20430] = 8'hf9 ;
            rom[20431] = 8'h12 ;
            rom[20432] = 8'hd0 ;
            rom[20433] = 8'he5 ;
            rom[20434] = 8'hec ;
            rom[20435] = 8'hfa ;
            rom[20436] = 8'h01 ;
            rom[20437] = 8'hf8 ;
            rom[20438] = 8'hea ;
            rom[20439] = 8'hf4 ;
            rom[20440] = 8'he4 ;
            rom[20441] = 8'hf1 ;
            rom[20442] = 8'hfa ;
            rom[20443] = 8'h14 ;
            rom[20444] = 8'ha7 ;
            rom[20445] = 8'h06 ;
            rom[20446] = 8'h11 ;
            rom[20447] = 8'h1d ;
            rom[20448] = 8'hfd ;
            rom[20449] = 8'hf2 ;
            rom[20450] = 8'h13 ;
            rom[20451] = 8'hfc ;
            rom[20452] = 8'hf6 ;
            rom[20453] = 8'hf0 ;
            rom[20454] = 8'h0b ;
            rom[20455] = 8'h07 ;
            rom[20456] = 8'hf3 ;
            rom[20457] = 8'hf8 ;
            rom[20458] = 8'hcd ;
            rom[20459] = 8'h18 ;
            rom[20460] = 8'hfc ;
            rom[20461] = 8'hfe ;
            rom[20462] = 8'h09 ;
            rom[20463] = 8'h0c ;
            rom[20464] = 8'he7 ;
            rom[20465] = 8'h04 ;
            rom[20466] = 8'he8 ;
            rom[20467] = 8'he0 ;
            rom[20468] = 8'hb3 ;
            rom[20469] = 8'h05 ;
            rom[20470] = 8'h06 ;
            rom[20471] = 8'hf6 ;
            rom[20472] = 8'hf9 ;
            rom[20473] = 8'h19 ;
            rom[20474] = 8'hec ;
            rom[20475] = 8'h05 ;
            rom[20476] = 8'hf7 ;
            rom[20477] = 8'he3 ;
            rom[20478] = 8'hed ;
            rom[20479] = 8'hf6 ;
            rom[20480] = 8'he0 ;
            rom[20481] = 8'hf6 ;
            rom[20482] = 8'hf7 ;
            rom[20483] = 8'h14 ;
            rom[20484] = 8'h05 ;
            rom[20485] = 8'hfc ;
            rom[20486] = 8'hfc ;
            rom[20487] = 8'h17 ;
            rom[20488] = 8'h26 ;
            rom[20489] = 8'he3 ;
            rom[20490] = 8'hf0 ;
            rom[20491] = 8'hf1 ;
            rom[20492] = 8'hfd ;
            rom[20493] = 8'h19 ;
            rom[20494] = 8'h0e ;
            rom[20495] = 8'hff ;
            rom[20496] = 8'hdd ;
            rom[20497] = 8'h1b ;
            rom[20498] = 8'h09 ;
            rom[20499] = 8'hbc ;
            rom[20500] = 8'hdc ;
            rom[20501] = 8'hf6 ;
            rom[20502] = 8'h18 ;
            rom[20503] = 8'h1d ;
            rom[20504] = 8'h06 ;
            rom[20505] = 8'h16 ;
            rom[20506] = 8'h04 ;
            rom[20507] = 8'he2 ;
            rom[20508] = 8'h02 ;
            rom[20509] = 8'hc9 ;
            rom[20510] = 8'h17 ;
            rom[20511] = 8'h02 ;
            rom[20512] = 8'he9 ;
            rom[20513] = 8'hd6 ;
            rom[20514] = 8'hf4 ;
            rom[20515] = 8'hc1 ;
            rom[20516] = 8'hdc ;
            rom[20517] = 8'hd8 ;
            rom[20518] = 8'h0d ;
            rom[20519] = 8'h12 ;
            rom[20520] = 8'hf7 ;
            rom[20521] = 8'hcc ;
            rom[20522] = 8'hf4 ;
            rom[20523] = 8'h13 ;
            rom[20524] = 8'h07 ;
            rom[20525] = 8'hcf ;
            rom[20526] = 8'h12 ;
            rom[20527] = 8'he3 ;
            rom[20528] = 8'h09 ;
            rom[20529] = 8'hfc ;
            rom[20530] = 8'hcc ;
            rom[20531] = 8'hde ;
            rom[20532] = 8'hea ;
            rom[20533] = 8'hd7 ;
            rom[20534] = 8'h19 ;
            rom[20535] = 8'hfd ;
            rom[20536] = 8'h09 ;
            rom[20537] = 8'hf3 ;
            rom[20538] = 8'hf8 ;
            rom[20539] = 8'hdb ;
            rom[20540] = 8'h12 ;
            rom[20541] = 8'hfa ;
            rom[20542] = 8'h02 ;
            rom[20543] = 8'h1a ;
            rom[20544] = 8'h1e ;
            rom[20545] = 8'he8 ;
            rom[20546] = 8'hf2 ;
            rom[20547] = 8'hce ;
            rom[20548] = 8'h0c ;
            rom[20549] = 8'hfd ;
            rom[20550] = 8'hf8 ;
            rom[20551] = 8'hff ;
            rom[20552] = 8'he4 ;
            rom[20553] = 8'hfe ;
            rom[20554] = 8'hc3 ;
            rom[20555] = 8'h04 ;
            rom[20556] = 8'hf4 ;
            rom[20557] = 8'h0f ;
            rom[20558] = 8'hd4 ;
            rom[20559] = 8'h15 ;
            rom[20560] = 8'h08 ;
            rom[20561] = 8'h1f ;
            rom[20562] = 8'h1d ;
            rom[20563] = 8'hde ;
            rom[20564] = 8'h1d ;
            rom[20565] = 8'he0 ;
            rom[20566] = 8'hef ;
            rom[20567] = 8'h19 ;
            rom[20568] = 8'hf1 ;
            rom[20569] = 8'hbe ;
            rom[20570] = 8'hea ;
            rom[20571] = 8'hf1 ;
            rom[20572] = 8'hf7 ;
            rom[20573] = 8'h23 ;
            rom[20574] = 8'hd0 ;
            rom[20575] = 8'hf1 ;
            rom[20576] = 8'h21 ;
            rom[20577] = 8'h0c ;
            rom[20578] = 8'he8 ;
            rom[20579] = 8'h05 ;
            rom[20580] = 8'h1a ;
            rom[20581] = 8'hff ;
            rom[20582] = 8'h20 ;
            rom[20583] = 8'h18 ;
            rom[20584] = 8'he5 ;
            rom[20585] = 8'h04 ;
            rom[20586] = 8'hdf ;
            rom[20587] = 8'h01 ;
            rom[20588] = 8'he7 ;
            rom[20589] = 8'h18 ;
            rom[20590] = 8'he9 ;
            rom[20591] = 8'he5 ;
            rom[20592] = 8'h31 ;
            rom[20593] = 8'h11 ;
            rom[20594] = 8'h17 ;
            rom[20595] = 8'h03 ;
            rom[20596] = 8'h18 ;
            rom[20597] = 8'h08 ;
            rom[20598] = 8'hd2 ;
            rom[20599] = 8'hbc ;
            rom[20600] = 8'hc9 ;
            rom[20601] = 8'h04 ;
            rom[20602] = 8'h07 ;
            rom[20603] = 8'h0d ;
            rom[20604] = 8'he3 ;
            rom[20605] = 8'he4 ;
            rom[20606] = 8'h02 ;
            rom[20607] = 8'h22 ;
            rom[20608] = 8'h29 ;
            rom[20609] = 8'hd7 ;
            rom[20610] = 8'hec ;
            rom[20611] = 8'h22 ;
            rom[20612] = 8'hff ;
            rom[20613] = 8'hff ;
            rom[20614] = 8'hf3 ;
            rom[20615] = 8'hd3 ;
            rom[20616] = 8'h13 ;
            rom[20617] = 8'h13 ;
            rom[20618] = 8'hfb ;
            rom[20619] = 8'hdd ;
            rom[20620] = 8'h02 ;
            rom[20621] = 8'he5 ;
            rom[20622] = 8'h16 ;
            rom[20623] = 8'h07 ;
            rom[20624] = 8'hea ;
            rom[20625] = 8'hf3 ;
            rom[20626] = 8'hf9 ;
            rom[20627] = 8'hf5 ;
            rom[20628] = 8'h02 ;
            rom[20629] = 8'he3 ;
            rom[20630] = 8'he1 ;
            rom[20631] = 8'h09 ;
            rom[20632] = 8'hfb ;
            rom[20633] = 8'hfc ;
            rom[20634] = 8'h03 ;
            rom[20635] = 8'hde ;
            rom[20636] = 8'hd8 ;
            rom[20637] = 8'h01 ;
            rom[20638] = 8'h0c ;
            rom[20639] = 8'h03 ;
            rom[20640] = 8'he4 ;
            rom[20641] = 8'hc9 ;
            rom[20642] = 8'hf9 ;
            rom[20643] = 8'hfe ;
            rom[20644] = 8'h12 ;
            rom[20645] = 8'h1e ;
            rom[20646] = 8'he3 ;
            rom[20647] = 8'hcf ;
            rom[20648] = 8'he8 ;
            rom[20649] = 8'hf4 ;
            rom[20650] = 8'h10 ;
            rom[20651] = 8'hf4 ;
            rom[20652] = 8'h05 ;
            rom[20653] = 8'h1c ;
            rom[20654] = 8'hec ;
            rom[20655] = 8'hea ;
            rom[20656] = 8'hf7 ;
            rom[20657] = 8'hf6 ;
            rom[20658] = 8'heb ;
            rom[20659] = 8'he4 ;
            rom[20660] = 8'hfe ;
            rom[20661] = 8'h01 ;
            rom[20662] = 8'heb ;
            rom[20663] = 8'hcf ;
            rom[20664] = 8'h0b ;
            rom[20665] = 8'hf3 ;
            rom[20666] = 8'h22 ;
            rom[20667] = 8'hf9 ;
            rom[20668] = 8'h1f ;
            rom[20669] = 8'hde ;
            rom[20670] = 8'h00 ;
            rom[20671] = 8'he3 ;
            rom[20672] = 8'hcf ;
            rom[20673] = 8'h22 ;
            rom[20674] = 8'hf5 ;
            rom[20675] = 8'h0c ;
            rom[20676] = 8'h19 ;
            rom[20677] = 8'hfb ;
            rom[20678] = 8'hdf ;
            rom[20679] = 8'h10 ;
            rom[20680] = 8'h1a ;
            rom[20681] = 8'hf7 ;
            rom[20682] = 8'hdd ;
            rom[20683] = 8'hf3 ;
            rom[20684] = 8'h28 ;
            rom[20685] = 8'h01 ;
            rom[20686] = 8'h33 ;
            rom[20687] = 8'h17 ;
            rom[20688] = 8'h28 ;
            rom[20689] = 8'hf9 ;
            rom[20690] = 8'hef ;
            rom[20691] = 8'hed ;
            rom[20692] = 8'he6 ;
            rom[20693] = 8'hfb ;
            rom[20694] = 8'hfb ;
            rom[20695] = 8'hfe ;
            rom[20696] = 8'h3d ;
            rom[20697] = 8'hd1 ;
            rom[20698] = 8'hfb ;
            rom[20699] = 8'h0c ;
            rom[20700] = 8'hf3 ;
            rom[20701] = 8'hfa ;
            rom[20702] = 8'hfa ;
            rom[20703] = 8'h12 ;
            rom[20704] = 8'hdc ;
            rom[20705] = 8'he6 ;
            rom[20706] = 8'h04 ;
            rom[20707] = 8'hff ;
            rom[20708] = 8'he4 ;
            rom[20709] = 8'hf6 ;
            rom[20710] = 8'h18 ;
            rom[20711] = 8'h0f ;
            rom[20712] = 8'hf5 ;
            rom[20713] = 8'hd8 ;
            rom[20714] = 8'hfe ;
            rom[20715] = 8'h29 ;
            rom[20716] = 8'h0a ;
            rom[20717] = 8'h08 ;
            rom[20718] = 8'h13 ;
            rom[20719] = 8'h10 ;
            rom[20720] = 8'hf9 ;
            rom[20721] = 8'hd8 ;
            rom[20722] = 8'h05 ;
            rom[20723] = 8'h09 ;
            rom[20724] = 8'h1f ;
            rom[20725] = 8'h1f ;
            rom[20726] = 8'h15 ;
            rom[20727] = 8'h12 ;
            rom[20728] = 8'h1e ;
            rom[20729] = 8'hf4 ;
            rom[20730] = 8'hd8 ;
            rom[20731] = 8'h01 ;
            rom[20732] = 8'he8 ;
            rom[20733] = 8'h03 ;
            rom[20734] = 8'hd2 ;
            rom[20735] = 8'hfe ;
            rom[20736] = 8'h00 ;
            rom[20737] = 8'h07 ;
            rom[20738] = 8'hf4 ;
            rom[20739] = 8'he8 ;
            rom[20740] = 8'h08 ;
            rom[20741] = 8'h08 ;
            rom[20742] = 8'he9 ;
            rom[20743] = 8'hea ;
            rom[20744] = 8'h06 ;
            rom[20745] = 8'h1d ;
            rom[20746] = 8'he2 ;
            rom[20747] = 8'hd3 ;
            rom[20748] = 8'h0b ;
            rom[20749] = 8'h04 ;
            rom[20750] = 8'h24 ;
            rom[20751] = 8'hf7 ;
            rom[20752] = 8'h18 ;
            rom[20753] = 8'h05 ;
            rom[20754] = 8'h0c ;
            rom[20755] = 8'hdb ;
            rom[20756] = 8'hf8 ;
            rom[20757] = 8'hf3 ;
            rom[20758] = 8'hf7 ;
            rom[20759] = 8'h07 ;
            rom[20760] = 8'hcc ;
            rom[20761] = 8'h03 ;
            rom[20762] = 8'hf0 ;
            rom[20763] = 8'heb ;
            rom[20764] = 8'hfb ;
            rom[20765] = 8'h03 ;
            rom[20766] = 8'h00 ;
            rom[20767] = 8'h04 ;
            rom[20768] = 8'h00 ;
            rom[20769] = 8'he7 ;
            rom[20770] = 8'hf6 ;
            rom[20771] = 8'he3 ;
            rom[20772] = 8'h13 ;
            rom[20773] = 8'hd6 ;
            rom[20774] = 8'h2c ;
            rom[20775] = 8'hea ;
            rom[20776] = 8'h01 ;
            rom[20777] = 8'hfd ;
            rom[20778] = 8'he8 ;
            rom[20779] = 8'hf3 ;
            rom[20780] = 8'hf7 ;
            rom[20781] = 8'hdd ;
            rom[20782] = 8'hf9 ;
            rom[20783] = 8'hfb ;
            rom[20784] = 8'h14 ;
            rom[20785] = 8'hfa ;
            rom[20786] = 8'heb ;
            rom[20787] = 8'h06 ;
            rom[20788] = 8'he9 ;
            rom[20789] = 8'hf3 ;
            rom[20790] = 8'h13 ;
            rom[20791] = 8'h06 ;
            rom[20792] = 8'hdd ;
            rom[20793] = 8'hc0 ;
            rom[20794] = 8'hf9 ;
            rom[20795] = 8'h27 ;
            rom[20796] = 8'h0e ;
            rom[20797] = 8'he7 ;
            rom[20798] = 8'h09 ;
            rom[20799] = 8'hff ;
            rom[20800] = 8'h07 ;
            rom[20801] = 8'hf1 ;
            rom[20802] = 8'h18 ;
            rom[20803] = 8'hf6 ;
            rom[20804] = 8'he2 ;
            rom[20805] = 8'hed ;
            rom[20806] = 8'h07 ;
            rom[20807] = 8'h08 ;
            rom[20808] = 8'h09 ;
            rom[20809] = 8'h01 ;
            rom[20810] = 8'hee ;
            rom[20811] = 8'h14 ;
            rom[20812] = 8'h0d ;
            rom[20813] = 8'hfd ;
            rom[20814] = 8'hde ;
            rom[20815] = 8'hd3 ;
            rom[20816] = 8'h00 ;
            rom[20817] = 8'h18 ;
            rom[20818] = 8'hf2 ;
            rom[20819] = 8'he5 ;
            rom[20820] = 8'hfc ;
            rom[20821] = 8'h1a ;
            rom[20822] = 8'hec ;
            rom[20823] = 8'h0c ;
            rom[20824] = 8'hf3 ;
            rom[20825] = 8'hbe ;
            rom[20826] = 8'hf5 ;
            rom[20827] = 8'h16 ;
            rom[20828] = 8'hd4 ;
            rom[20829] = 8'h04 ;
            rom[20830] = 8'hde ;
            rom[20831] = 8'hfe ;
            rom[20832] = 8'hd6 ;
            rom[20833] = 8'h0c ;
            rom[20834] = 8'h0f ;
            rom[20835] = 8'hf9 ;
            rom[20836] = 8'h08 ;
            rom[20837] = 8'h04 ;
            rom[20838] = 8'h11 ;
            rom[20839] = 8'hf2 ;
            rom[20840] = 8'hf7 ;
            rom[20841] = 8'hed ;
            rom[20842] = 8'h30 ;
            rom[20843] = 8'h2b ;
            rom[20844] = 8'h2c ;
            rom[20845] = 8'hd0 ;
            rom[20846] = 8'hec ;
            rom[20847] = 8'hfb ;
            rom[20848] = 8'h01 ;
            rom[20849] = 8'h16 ;
            rom[20850] = 8'h07 ;
            rom[20851] = 8'h0d ;
            rom[20852] = 8'h25 ;
            rom[20853] = 8'hf2 ;
            rom[20854] = 8'hda ;
            rom[20855] = 8'h07 ;
            rom[20856] = 8'h10 ;
            rom[20857] = 8'h1c ;
            rom[20858] = 8'hfa ;
            rom[20859] = 8'hf7 ;
            rom[20860] = 8'h19 ;
            rom[20861] = 8'h21 ;
            rom[20862] = 8'hf7 ;
            rom[20863] = 8'hec ;
            rom[20864] = 8'h0e ;
            rom[20865] = 8'hce ;
            rom[20866] = 8'hf4 ;
            rom[20867] = 8'hff ;
            rom[20868] = 8'he4 ;
            rom[20869] = 8'h05 ;
            rom[20870] = 8'hee ;
            rom[20871] = 8'hee ;
            rom[20872] = 8'h08 ;
            rom[20873] = 8'h12 ;
            rom[20874] = 8'h01 ;
            rom[20875] = 8'h19 ;
            rom[20876] = 8'h11 ;
            rom[20877] = 8'hea ;
            rom[20878] = 8'h15 ;
            rom[20879] = 8'hf9 ;
            rom[20880] = 8'hc1 ;
            rom[20881] = 8'hcc ;
            rom[20882] = 8'h13 ;
            rom[20883] = 8'h08 ;
            rom[20884] = 8'h10 ;
            rom[20885] = 8'hed ;
            rom[20886] = 8'hed ;
            rom[20887] = 8'h1f ;
            rom[20888] = 8'hec ;
            rom[20889] = 8'h0e ;
            rom[20890] = 8'h20 ;
            rom[20891] = 8'hbb ;
            rom[20892] = 8'hde ;
            rom[20893] = 8'he3 ;
            rom[20894] = 8'h09 ;
            rom[20895] = 8'h24 ;
            rom[20896] = 8'hfb ;
            rom[20897] = 8'hcf ;
            rom[20898] = 8'hf2 ;
            rom[20899] = 8'h1b ;
            rom[20900] = 8'h1f ;
            rom[20901] = 8'h09 ;
            rom[20902] = 8'h0b ;
            rom[20903] = 8'he9 ;
            rom[20904] = 8'h05 ;
            rom[20905] = 8'hd5 ;
            rom[20906] = 8'hf4 ;
            rom[20907] = 8'hfd ;
            rom[20908] = 8'hf0 ;
            rom[20909] = 8'h19 ;
            rom[20910] = 8'he0 ;
            rom[20911] = 8'hf5 ;
            rom[20912] = 8'he5 ;
            rom[20913] = 8'hdc ;
            rom[20914] = 8'h0b ;
            rom[20915] = 8'hd2 ;
            rom[20916] = 8'hf0 ;
            rom[20917] = 8'h05 ;
            rom[20918] = 8'hea ;
            rom[20919] = 8'ha3 ;
            rom[20920] = 8'hff ;
            rom[20921] = 8'hd7 ;
            rom[20922] = 8'h02 ;
            rom[20923] = 8'h10 ;
            rom[20924] = 8'h09 ;
            rom[20925] = 8'hfc ;
            rom[20926] = 8'hf9 ;
            rom[20927] = 8'hea ;
            rom[20928] = 8'hd9 ;
            rom[20929] = 8'h16 ;
            rom[20930] = 8'h20 ;
            rom[20931] = 8'hf4 ;
            rom[20932] = 8'h06 ;
            rom[20933] = 8'h01 ;
            rom[20934] = 8'hf3 ;
            rom[20935] = 8'h20 ;
            rom[20936] = 8'h13 ;
            rom[20937] = 8'h14 ;
            rom[20938] = 8'hd1 ;
            rom[20939] = 8'he7 ;
            rom[20940] = 8'hec ;
            rom[20941] = 8'h17 ;
            rom[20942] = 8'h2c ;
            rom[20943] = 8'he3 ;
            rom[20944] = 8'h1f ;
            rom[20945] = 8'hfb ;
            rom[20946] = 8'he6 ;
            rom[20947] = 8'he7 ;
            rom[20948] = 8'hf1 ;
            rom[20949] = 8'he8 ;
            rom[20950] = 8'h17 ;
            rom[20951] = 8'hc5 ;
            rom[20952] = 8'h04 ;
            rom[20953] = 8'hd6 ;
            rom[20954] = 8'hfc ;
            rom[20955] = 8'h20 ;
            rom[20956] = 8'hf0 ;
            rom[20957] = 8'hf4 ;
            rom[20958] = 8'h06 ;
            rom[20959] = 8'h02 ;
            rom[20960] = 8'hd3 ;
            rom[20961] = 8'h00 ;
            rom[20962] = 8'hf0 ;
            rom[20963] = 8'hf7 ;
            rom[20964] = 8'hfd ;
            rom[20965] = 8'hf6 ;
            rom[20966] = 8'h0a ;
            rom[20967] = 8'hfd ;
            rom[20968] = 8'hdf ;
            rom[20969] = 8'hc3 ;
            rom[20970] = 8'h13 ;
            rom[20971] = 8'hf4 ;
            rom[20972] = 8'h0b ;
            rom[20973] = 8'h14 ;
            rom[20974] = 8'h0f ;
            rom[20975] = 8'hfd ;
            rom[20976] = 8'hf6 ;
            rom[20977] = 8'h09 ;
            rom[20978] = 8'h29 ;
            rom[20979] = 8'h0c ;
            rom[20980] = 8'h1f ;
            rom[20981] = 8'h1d ;
            rom[20982] = 8'hfc ;
            rom[20983] = 8'hcd ;
            rom[20984] = 8'hfe ;
            rom[20985] = 8'h03 ;
            rom[20986] = 8'he8 ;
            rom[20987] = 8'hc8 ;
            rom[20988] = 8'hf6 ;
            rom[20989] = 8'h0f ;
            rom[20990] = 8'hd7 ;
            rom[20991] = 8'hfa ;
            rom[20992] = 8'h06 ;
            rom[20993] = 8'h11 ;
            rom[20994] = 8'hf0 ;
            rom[20995] = 8'he3 ;
            rom[20996] = 8'h18 ;
            rom[20997] = 8'h09 ;
            rom[20998] = 8'hfa ;
            rom[20999] = 8'hfa ;
            rom[21000] = 8'he8 ;
            rom[21001] = 8'he3 ;
            rom[21002] = 8'h01 ;
            rom[21003] = 8'h0b ;
            rom[21004] = 8'h0a ;
            rom[21005] = 8'he3 ;
            rom[21006] = 8'hc6 ;
            rom[21007] = 8'hfa ;
            rom[21008] = 8'hf6 ;
            rom[21009] = 8'heb ;
            rom[21010] = 8'h1e ;
            rom[21011] = 8'hea ;
            rom[21012] = 8'h1b ;
            rom[21013] = 8'h05 ;
            rom[21014] = 8'hfa ;
            rom[21015] = 8'hfc ;
            rom[21016] = 8'h28 ;
            rom[21017] = 8'h0b ;
            rom[21018] = 8'heb ;
            rom[21019] = 8'hed ;
            rom[21020] = 8'h04 ;
            rom[21021] = 8'h24 ;
            rom[21022] = 8'hec ;
            rom[21023] = 8'h15 ;
            rom[21024] = 8'h0e ;
            rom[21025] = 8'h02 ;
            rom[21026] = 8'h01 ;
            rom[21027] = 8'h00 ;
            rom[21028] = 8'h06 ;
            rom[21029] = 8'hdb ;
            rom[21030] = 8'hf7 ;
            rom[21031] = 8'hdb ;
            rom[21032] = 8'h38 ;
            rom[21033] = 8'he5 ;
            rom[21034] = 8'hdd ;
            rom[21035] = 8'hf5 ;
            rom[21036] = 8'hf6 ;
            rom[21037] = 8'h1f ;
            rom[21038] = 8'he9 ;
            rom[21039] = 8'he4 ;
            rom[21040] = 8'hef ;
            rom[21041] = 8'h26 ;
            rom[21042] = 8'h06 ;
            rom[21043] = 8'hff ;
            rom[21044] = 8'h0b ;
            rom[21045] = 8'hff ;
            rom[21046] = 8'hef ;
            rom[21047] = 8'hfb ;
            rom[21048] = 8'hf3 ;
            rom[21049] = 8'h12 ;
            rom[21050] = 8'hd4 ;
            rom[21051] = 8'he9 ;
            rom[21052] = 8'hf2 ;
            rom[21053] = 8'hd7 ;
            rom[21054] = 8'hc2 ;
            rom[21055] = 8'h01 ;
            rom[21056] = 8'hff ;
            rom[21057] = 8'h18 ;
            rom[21058] = 8'h0d ;
            rom[21059] = 8'h14 ;
            rom[21060] = 8'h03 ;
            rom[21061] = 8'h0e ;
            rom[21062] = 8'he8 ;
            rom[21063] = 8'h02 ;
            rom[21064] = 8'hd4 ;
            rom[21065] = 8'h02 ;
            rom[21066] = 8'h01 ;
            rom[21067] = 8'hf7 ;
            rom[21068] = 8'hf6 ;
            rom[21069] = 8'he0 ;
            rom[21070] = 8'heb ;
            rom[21071] = 8'h0a ;
            rom[21072] = 8'h00 ;
            rom[21073] = 8'hf2 ;
            rom[21074] = 8'h1b ;
            rom[21075] = 8'h0e ;
            rom[21076] = 8'hb0 ;
            rom[21077] = 8'h04 ;
            rom[21078] = 8'h0f ;
            rom[21079] = 8'hee ;
            rom[21080] = 8'hf7 ;
            rom[21081] = 8'hf1 ;
            rom[21082] = 8'h1f ;
            rom[21083] = 8'h29 ;
            rom[21084] = 8'h03 ;
            rom[21085] = 8'h0c ;
            rom[21086] = 8'hf1 ;
            rom[21087] = 8'hef ;
            rom[21088] = 8'h0f ;
            rom[21089] = 8'h0b ;
            rom[21090] = 8'h03 ;
            rom[21091] = 8'hfd ;
            rom[21092] = 8'h09 ;
            rom[21093] = 8'h44 ;
            rom[21094] = 8'h14 ;
            rom[21095] = 8'hf0 ;
            rom[21096] = 8'h0d ;
            rom[21097] = 8'hf5 ;
            rom[21098] = 8'hfc ;
            rom[21099] = 8'h2f ;
            rom[21100] = 8'hec ;
            rom[21101] = 8'hfb ;
            rom[21102] = 8'he2 ;
            rom[21103] = 8'h1d ;
            rom[21104] = 8'hf8 ;
            rom[21105] = 8'he8 ;
            rom[21106] = 8'hdd ;
            rom[21107] = 8'h0a ;
            rom[21108] = 8'hc9 ;
            rom[21109] = 8'h0a ;
            rom[21110] = 8'hed ;
            rom[21111] = 8'he8 ;
            rom[21112] = 8'hdf ;
            rom[21113] = 8'h0c ;
            rom[21114] = 8'hf9 ;
            rom[21115] = 8'he2 ;
            rom[21116] = 8'h11 ;
            rom[21117] = 8'h0f ;
            rom[21118] = 8'h01 ;
            rom[21119] = 8'h1f ;
            rom[21120] = 8'he6 ;
            rom[21121] = 8'h17 ;
            rom[21122] = 8'hfd ;
            rom[21123] = 8'hf7 ;
            rom[21124] = 8'h08 ;
            rom[21125] = 8'h03 ;
            rom[21126] = 8'h18 ;
            rom[21127] = 8'hf0 ;
            rom[21128] = 8'h03 ;
            rom[21129] = 8'he0 ;
            rom[21130] = 8'h0f ;
            rom[21131] = 8'hfc ;
            rom[21132] = 8'hef ;
            rom[21133] = 8'hfb ;
            rom[21134] = 8'he1 ;
            rom[21135] = 8'h0a ;
            rom[21136] = 8'h19 ;
            rom[21137] = 8'h24 ;
            rom[21138] = 8'he2 ;
            rom[21139] = 8'hcc ;
            rom[21140] = 8'h0a ;
            rom[21141] = 8'h05 ;
            rom[21142] = 8'he2 ;
            rom[21143] = 8'hdf ;
            rom[21144] = 8'hfc ;
            rom[21145] = 8'hef ;
            rom[21146] = 8'h10 ;
            rom[21147] = 8'h26 ;
            rom[21148] = 8'h25 ;
            rom[21149] = 8'h20 ;
            rom[21150] = 8'hd7 ;
            rom[21151] = 8'hd6 ;
            rom[21152] = 8'h2b ;
            rom[21153] = 8'h0f ;
            rom[21154] = 8'h23 ;
            rom[21155] = 8'h02 ;
            rom[21156] = 8'he0 ;
            rom[21157] = 8'h12 ;
            rom[21158] = 8'he7 ;
            rom[21159] = 8'h18 ;
            rom[21160] = 8'h00 ;
            rom[21161] = 8'h04 ;
            rom[21162] = 8'hf9 ;
            rom[21163] = 8'hfc ;
            rom[21164] = 8'h13 ;
            rom[21165] = 8'h0b ;
            rom[21166] = 8'h18 ;
            rom[21167] = 8'hea ;
            rom[21168] = 8'hf0 ;
            rom[21169] = 8'hf3 ;
            rom[21170] = 8'hef ;
            rom[21171] = 8'he1 ;
            rom[21172] = 8'h01 ;
            rom[21173] = 8'hf6 ;
            rom[21174] = 8'h00 ;
            rom[21175] = 8'h15 ;
            rom[21176] = 8'h21 ;
            rom[21177] = 8'hee ;
            rom[21178] = 8'he5 ;
            rom[21179] = 8'hca ;
            rom[21180] = 8'hf8 ;
            rom[21181] = 8'he2 ;
            rom[21182] = 8'hff ;
            rom[21183] = 8'hf0 ;
            rom[21184] = 8'hf2 ;
            rom[21185] = 8'hed ;
            rom[21186] = 8'hec ;
            rom[21187] = 8'h19 ;
            rom[21188] = 8'hfe ;
            rom[21189] = 8'hfc ;
            rom[21190] = 8'hf4 ;
            rom[21191] = 8'h28 ;
            rom[21192] = 8'hd2 ;
            rom[21193] = 8'h04 ;
            rom[21194] = 8'hfb ;
            rom[21195] = 8'h26 ;
            rom[21196] = 8'hf5 ;
            rom[21197] = 8'he7 ;
            rom[21198] = 8'hf6 ;
            rom[21199] = 8'hf2 ;
            rom[21200] = 8'h0d ;
            rom[21201] = 8'hd3 ;
            rom[21202] = 8'hf7 ;
            rom[21203] = 8'hfd ;
            rom[21204] = 8'h0c ;
            rom[21205] = 8'hfc ;
            rom[21206] = 8'h03 ;
            rom[21207] = 8'hee ;
            rom[21208] = 8'hf8 ;
            rom[21209] = 8'hf5 ;
            rom[21210] = 8'h11 ;
            rom[21211] = 8'h11 ;
            rom[21212] = 8'h38 ;
            rom[21213] = 8'h19 ;
            rom[21214] = 8'h18 ;
            rom[21215] = 8'h05 ;
            rom[21216] = 8'he6 ;
            rom[21217] = 8'hef ;
            rom[21218] = 8'h23 ;
            rom[21219] = 8'he5 ;
            rom[21220] = 8'h02 ;
            rom[21221] = 8'h05 ;
            rom[21222] = 8'h19 ;
            rom[21223] = 8'hfd ;
            rom[21224] = 8'h08 ;
            rom[21225] = 8'h1e ;
            rom[21226] = 8'h1c ;
            rom[21227] = 8'hf4 ;
            rom[21228] = 8'h1c ;
            rom[21229] = 8'hde ;
            rom[21230] = 8'hf9 ;
            rom[21231] = 8'h08 ;
            rom[21232] = 8'h06 ;
            rom[21233] = 8'hfb ;
            rom[21234] = 8'h34 ;
            rom[21235] = 8'h16 ;
            rom[21236] = 8'h0d ;
            rom[21237] = 8'h0e ;
            rom[21238] = 8'he6 ;
            rom[21239] = 8'h00 ;
            rom[21240] = 8'he7 ;
            rom[21241] = 8'hcf ;
            rom[21242] = 8'hf3 ;
            rom[21243] = 8'hf1 ;
            rom[21244] = 8'h02 ;
            rom[21245] = 8'h17 ;
            rom[21246] = 8'hfb ;
            rom[21247] = 8'h13 ;
            rom[21248] = 8'hcc ;
            rom[21249] = 8'he4 ;
            rom[21250] = 8'h0e ;
            rom[21251] = 8'h17 ;
            rom[21252] = 8'hdd ;
            rom[21253] = 8'hfd ;
            rom[21254] = 8'h0c ;
            rom[21255] = 8'hf2 ;
            rom[21256] = 8'h1d ;
            rom[21257] = 8'hfe ;
            rom[21258] = 8'h00 ;
            rom[21259] = 8'he8 ;
            rom[21260] = 8'h27 ;
            rom[21261] = 8'hd9 ;
            rom[21262] = 8'h2b ;
            rom[21263] = 8'h0e ;
            rom[21264] = 8'hc0 ;
            rom[21265] = 8'h01 ;
            rom[21266] = 8'h0a ;
            rom[21267] = 8'h07 ;
            rom[21268] = 8'hf1 ;
            rom[21269] = 8'he3 ;
            rom[21270] = 8'hee ;
            rom[21271] = 8'h2c ;
            rom[21272] = 8'hfa ;
            rom[21273] = 8'h30 ;
            rom[21274] = 8'h2d ;
            rom[21275] = 8'h10 ;
            rom[21276] = 8'h09 ;
            rom[21277] = 8'hd8 ;
            rom[21278] = 8'h0e ;
            rom[21279] = 8'he7 ;
            rom[21280] = 8'hfa ;
            rom[21281] = 8'hb5 ;
            rom[21282] = 8'he7 ;
            rom[21283] = 8'hf7 ;
            rom[21284] = 8'h00 ;
            rom[21285] = 8'h0d ;
            rom[21286] = 8'hff ;
            rom[21287] = 8'hfa ;
            rom[21288] = 8'h14 ;
            rom[21289] = 8'hbe ;
            rom[21290] = 8'hf3 ;
            rom[21291] = 8'hf0 ;
            rom[21292] = 8'hd8 ;
            rom[21293] = 8'he6 ;
            rom[21294] = 8'hd3 ;
            rom[21295] = 8'hee ;
            rom[21296] = 8'he7 ;
            rom[21297] = 8'h24 ;
            rom[21298] = 8'hf6 ;
            rom[21299] = 8'hf9 ;
            rom[21300] = 8'h06 ;
            rom[21301] = 8'hf9 ;
            rom[21302] = 8'hd1 ;
            rom[21303] = 8'h02 ;
            rom[21304] = 8'he0 ;
            rom[21305] = 8'h06 ;
            rom[21306] = 8'h1e ;
            rom[21307] = 8'he8 ;
            rom[21308] = 8'h11 ;
            rom[21309] = 8'h01 ;
            rom[21310] = 8'hfb ;
            rom[21311] = 8'hf8 ;
            rom[21312] = 8'hc7 ;
            rom[21313] = 8'hf9 ;
            rom[21314] = 8'h02 ;
            rom[21315] = 8'hfe ;
            rom[21316] = 8'hf1 ;
            rom[21317] = 8'h0b ;
            rom[21318] = 8'hf3 ;
            rom[21319] = 8'h00 ;
            rom[21320] = 8'h27 ;
            rom[21321] = 8'h0c ;
            rom[21322] = 8'he6 ;
            rom[21323] = 8'h00 ;
            rom[21324] = 8'h27 ;
            rom[21325] = 8'h24 ;
            rom[21326] = 8'h1b ;
            rom[21327] = 8'hdb ;
            rom[21328] = 8'hf2 ;
            rom[21329] = 8'hea ;
            rom[21330] = 8'h05 ;
            rom[21331] = 8'hec ;
            rom[21332] = 8'h03 ;
            rom[21333] = 8'hef ;
            rom[21334] = 8'h0e ;
            rom[21335] = 8'h10 ;
            rom[21336] = 8'h0f ;
            rom[21337] = 8'he5 ;
            rom[21338] = 8'h01 ;
            rom[21339] = 8'h11 ;
            rom[21340] = 8'h1a ;
            rom[21341] = 8'hee ;
            rom[21342] = 8'h0e ;
            rom[21343] = 8'h0b ;
            rom[21344] = 8'hfa ;
            rom[21345] = 8'h01 ;
            rom[21346] = 8'hf8 ;
            rom[21347] = 8'h3c ;
            rom[21348] = 8'h1c ;
            rom[21349] = 8'h16 ;
            rom[21350] = 8'h2c ;
            rom[21351] = 8'h0e ;
            rom[21352] = 8'hf4 ;
            rom[21353] = 8'h0d ;
            rom[21354] = 8'hef ;
            rom[21355] = 8'hff ;
            rom[21356] = 8'h00 ;
            rom[21357] = 8'h0c ;
            rom[21358] = 8'hf6 ;
            rom[21359] = 8'hc4 ;
            rom[21360] = 8'h00 ;
            rom[21361] = 8'h03 ;
            rom[21362] = 8'hf1 ;
            rom[21363] = 8'hec ;
            rom[21364] = 8'h0f ;
            rom[21365] = 8'h01 ;
            rom[21366] = 8'hf8 ;
            rom[21367] = 8'he4 ;
            rom[21368] = 8'hf0 ;
            rom[21369] = 8'h04 ;
            rom[21370] = 8'h37 ;
            rom[21371] = 8'h0b ;
            rom[21372] = 8'hce ;
            rom[21373] = 8'heb ;
            rom[21374] = 8'hff ;
            rom[21375] = 8'h10 ;
            rom[21376] = 8'h02 ;
            rom[21377] = 8'he9 ;
            rom[21378] = 8'hf5 ;
            rom[21379] = 8'he0 ;
            rom[21380] = 8'heb ;
            rom[21381] = 8'h0a ;
            rom[21382] = 8'h08 ;
            rom[21383] = 8'hf0 ;
            rom[21384] = 8'hfa ;
            rom[21385] = 8'h08 ;
            rom[21386] = 8'hd9 ;
            rom[21387] = 8'h14 ;
            rom[21388] = 8'hfe ;
            rom[21389] = 8'h04 ;
            rom[21390] = 8'h0b ;
            rom[21391] = 8'h07 ;
            rom[21392] = 8'h26 ;
            rom[21393] = 8'h0e ;
            rom[21394] = 8'h01 ;
            rom[21395] = 8'h03 ;
            rom[21396] = 8'h3e ;
            rom[21397] = 8'h02 ;
            rom[21398] = 8'h00 ;
            rom[21399] = 8'hfe ;
            rom[21400] = 8'hd6 ;
            rom[21401] = 8'h12 ;
            rom[21402] = 8'h1a ;
            rom[21403] = 8'hef ;
            rom[21404] = 8'hf5 ;
            rom[21405] = 8'h04 ;
            rom[21406] = 8'h0a ;
            rom[21407] = 8'h1b ;
            rom[21408] = 8'heb ;
            rom[21409] = 8'hf3 ;
            rom[21410] = 8'h1a ;
            rom[21411] = 8'hd7 ;
            rom[21412] = 8'hf3 ;
            rom[21413] = 8'h0d ;
            rom[21414] = 8'hfe ;
            rom[21415] = 8'hed ;
            rom[21416] = 8'hf3 ;
            rom[21417] = 8'h08 ;
            rom[21418] = 8'h11 ;
            rom[21419] = 8'h23 ;
            rom[21420] = 8'hfc ;
            rom[21421] = 8'hfb ;
            rom[21422] = 8'hf6 ;
            rom[21423] = 8'hf2 ;
            rom[21424] = 8'h09 ;
            rom[21425] = 8'he4 ;
            rom[21426] = 8'h21 ;
            rom[21427] = 8'hdf ;
            rom[21428] = 8'hf5 ;
            rom[21429] = 8'hf9 ;
            rom[21430] = 8'h07 ;
            rom[21431] = 8'hd8 ;
            rom[21432] = 8'hf7 ;
            rom[21433] = 8'he6 ;
            rom[21434] = 8'h0c ;
            rom[21435] = 8'h0f ;
            rom[21436] = 8'hf0 ;
            rom[21437] = 8'hd2 ;
            rom[21438] = 8'h0d ;
            rom[21439] = 8'h16 ;
            rom[21440] = 8'hcd ;
            rom[21441] = 8'hf1 ;
            rom[21442] = 8'h15 ;
            rom[21443] = 8'hf1 ;
            rom[21444] = 8'h11 ;
            rom[21445] = 8'h0d ;
            rom[21446] = 8'h18 ;
            rom[21447] = 8'hf9 ;
            rom[21448] = 8'h12 ;
            rom[21449] = 8'h05 ;
            rom[21450] = 8'hf1 ;
            rom[21451] = 8'hfc ;
            rom[21452] = 8'h02 ;
            rom[21453] = 8'hda ;
            rom[21454] = 8'hff ;
            rom[21455] = 8'hf8 ;
            rom[21456] = 8'hed ;
            rom[21457] = 8'hfb ;
            rom[21458] = 8'he7 ;
            rom[21459] = 8'he1 ;
            rom[21460] = 8'h0c ;
            rom[21461] = 8'hea ;
            rom[21462] = 8'he3 ;
            rom[21463] = 8'h2a ;
            rom[21464] = 8'h07 ;
            rom[21465] = 8'hd8 ;
            rom[21466] = 8'h03 ;
            rom[21467] = 8'h0e ;
            rom[21468] = 8'h03 ;
            rom[21469] = 8'he7 ;
            rom[21470] = 8'h09 ;
            rom[21471] = 8'h15 ;
            rom[21472] = 8'hf9 ;
            rom[21473] = 8'h04 ;
            rom[21474] = 8'h00 ;
            rom[21475] = 8'hd6 ;
            rom[21476] = 8'heb ;
            rom[21477] = 8'h11 ;
            rom[21478] = 8'hdb ;
            rom[21479] = 8'h03 ;
            rom[21480] = 8'hee ;
            rom[21481] = 8'h08 ;
            rom[21482] = 8'h1a ;
            rom[21483] = 8'he6 ;
            rom[21484] = 8'h16 ;
            rom[21485] = 8'h10 ;
            rom[21486] = 8'h01 ;
            rom[21487] = 8'hec ;
            rom[21488] = 8'he8 ;
            rom[21489] = 8'h0a ;
            rom[21490] = 8'h04 ;
            rom[21491] = 8'hf7 ;
            rom[21492] = 8'hdd ;
            rom[21493] = 8'he9 ;
            rom[21494] = 8'hed ;
            rom[21495] = 8'h14 ;
            rom[21496] = 8'h3b ;
            rom[21497] = 8'hd9 ;
            rom[21498] = 8'hd1 ;
            rom[21499] = 8'hda ;
            rom[21500] = 8'hfe ;
            rom[21501] = 8'h0e ;
            rom[21502] = 8'hed ;
            rom[21503] = 8'hda ;
            rom[21504] = 8'h02 ;
            rom[21505] = 8'hfa ;
            rom[21506] = 8'hff ;
            rom[21507] = 8'h0e ;
            rom[21508] = 8'h17 ;
            rom[21509] = 8'he4 ;
            rom[21510] = 8'h0e ;
            rom[21511] = 8'h02 ;
            rom[21512] = 8'h00 ;
            rom[21513] = 8'hed ;
            rom[21514] = 8'h1e ;
            rom[21515] = 8'hef ;
            rom[21516] = 8'h1a ;
            rom[21517] = 8'hf1 ;
            rom[21518] = 8'hfe ;
            rom[21519] = 8'hdd ;
            rom[21520] = 8'hcf ;
            rom[21521] = 8'hfc ;
            rom[21522] = 8'h42 ;
            rom[21523] = 8'hc8 ;
            rom[21524] = 8'hdb ;
            rom[21525] = 8'hf2 ;
            rom[21526] = 8'h17 ;
            rom[21527] = 8'hed ;
            rom[21528] = 8'hd2 ;
            rom[21529] = 8'h1d ;
            rom[21530] = 8'h03 ;
            rom[21531] = 8'hea ;
            rom[21532] = 8'h03 ;
            rom[21533] = 8'hff ;
            rom[21534] = 8'h07 ;
            rom[21535] = 8'hfa ;
            rom[21536] = 8'heb ;
            rom[21537] = 8'h13 ;
            rom[21538] = 8'hf7 ;
            rom[21539] = 8'h01 ;
            rom[21540] = 8'he4 ;
            rom[21541] = 8'h07 ;
            rom[21542] = 8'h1a ;
            rom[21543] = 8'he1 ;
            rom[21544] = 8'hf8 ;
            rom[21545] = 8'h00 ;
            rom[21546] = 8'hff ;
            rom[21547] = 8'h09 ;
            rom[21548] = 8'hf9 ;
            rom[21549] = 8'hf4 ;
            rom[21550] = 8'h09 ;
            rom[21551] = 8'h02 ;
            rom[21552] = 8'h19 ;
            rom[21553] = 8'he5 ;
            rom[21554] = 8'he6 ;
            rom[21555] = 8'h05 ;
            rom[21556] = 8'hee ;
            rom[21557] = 8'hf1 ;
            rom[21558] = 8'h08 ;
            rom[21559] = 8'hf7 ;
            rom[21560] = 8'h03 ;
            rom[21561] = 8'hf4 ;
            rom[21562] = 8'h03 ;
            rom[21563] = 8'he1 ;
            rom[21564] = 8'h02 ;
            rom[21565] = 8'h0b ;
            rom[21566] = 8'h08 ;
            rom[21567] = 8'h0a ;
            rom[21568] = 8'h06 ;
            rom[21569] = 8'hf0 ;
            rom[21570] = 8'hf9 ;
            rom[21571] = 8'he9 ;
            rom[21572] = 8'hfd ;
            rom[21573] = 8'h06 ;
            rom[21574] = 8'h08 ;
            rom[21575] = 8'hf5 ;
            rom[21576] = 8'heb ;
            rom[21577] = 8'hbe ;
            rom[21578] = 8'h03 ;
            rom[21579] = 8'hfc ;
            rom[21580] = 8'hf0 ;
            rom[21581] = 8'h03 ;
            rom[21582] = 8'hbc ;
            rom[21583] = 8'hf6 ;
            rom[21584] = 8'h14 ;
            rom[21585] = 8'h04 ;
            rom[21586] = 8'h04 ;
            rom[21587] = 8'h0a ;
            rom[21588] = 8'h1f ;
            rom[21589] = 8'hea ;
            rom[21590] = 8'hea ;
            rom[21591] = 8'h0a ;
            rom[21592] = 8'he4 ;
            rom[21593] = 8'hec ;
            rom[21594] = 8'hf2 ;
            rom[21595] = 8'hf1 ;
            rom[21596] = 8'hde ;
            rom[21597] = 8'hff ;
            rom[21598] = 8'h03 ;
            rom[21599] = 8'h04 ;
            rom[21600] = 8'h00 ;
            rom[21601] = 8'h00 ;
            rom[21602] = 8'hb6 ;
            rom[21603] = 8'h13 ;
            rom[21604] = 8'h1d ;
            rom[21605] = 8'hfd ;
            rom[21606] = 8'h28 ;
            rom[21607] = 8'h09 ;
            rom[21608] = 8'hcb ;
            rom[21609] = 8'hf3 ;
            rom[21610] = 8'hde ;
            rom[21611] = 8'hf9 ;
            rom[21612] = 8'hdd ;
            rom[21613] = 8'h1a ;
            rom[21614] = 8'hf3 ;
            rom[21615] = 8'h0b ;
            rom[21616] = 8'he6 ;
            rom[21617] = 8'h0f ;
            rom[21618] = 8'h3a ;
            rom[21619] = 8'hfe ;
            rom[21620] = 8'hde ;
            rom[21621] = 8'he7 ;
            rom[21622] = 8'hfa ;
            rom[21623] = 8'hc9 ;
            rom[21624] = 8'hdc ;
            rom[21625] = 8'h00 ;
            rom[21626] = 8'hf6 ;
            rom[21627] = 8'h1d ;
            rom[21628] = 8'h15 ;
            rom[21629] = 8'he6 ;
            rom[21630] = 8'h32 ;
            rom[21631] = 8'hff ;
            rom[21632] = 8'h1d ;
            rom[21633] = 8'hd0 ;
            rom[21634] = 8'he5 ;
            rom[21635] = 8'h00 ;
            rom[21636] = 8'hdf ;
            rom[21637] = 8'hd7 ;
            rom[21638] = 8'hf9 ;
            rom[21639] = 8'hfe ;
            rom[21640] = 8'hff ;
            rom[21641] = 8'hfc ;
            rom[21642] = 8'hf5 ;
            rom[21643] = 8'hef ;
            rom[21644] = 8'hf4 ;
            rom[21645] = 8'hea ;
            rom[21646] = 8'hda ;
            rom[21647] = 8'he3 ;
            rom[21648] = 8'h00 ;
            rom[21649] = 8'hf0 ;
            rom[21650] = 8'hfc ;
            rom[21651] = 8'h13 ;
            rom[21652] = 8'h13 ;
            rom[21653] = 8'hed ;
            rom[21654] = 8'hca ;
            rom[21655] = 8'h06 ;
            rom[21656] = 8'hcf ;
            rom[21657] = 8'h1c ;
            rom[21658] = 8'h18 ;
            rom[21659] = 8'hed ;
            rom[21660] = 8'hfb ;
            rom[21661] = 8'h03 ;
            rom[21662] = 8'hfe ;
            rom[21663] = 8'h06 ;
            rom[21664] = 8'h16 ;
            rom[21665] = 8'h0b ;
            rom[21666] = 8'h02 ;
            rom[21667] = 8'h09 ;
            rom[21668] = 8'h0b ;
            rom[21669] = 8'hde ;
            rom[21670] = 8'hca ;
            rom[21671] = 8'he0 ;
            rom[21672] = 8'hd0 ;
            rom[21673] = 8'h0e ;
            rom[21674] = 8'h12 ;
            rom[21675] = 8'hf6 ;
            rom[21676] = 8'hf5 ;
            rom[21677] = 8'h07 ;
            rom[21678] = 8'he0 ;
            rom[21679] = 8'h15 ;
            rom[21680] = 8'hfb ;
            rom[21681] = 8'he9 ;
            rom[21682] = 8'h05 ;
            rom[21683] = 8'heb ;
            rom[21684] = 8'h13 ;
            rom[21685] = 8'h0e ;
            rom[21686] = 8'hca ;
            rom[21687] = 8'hea ;
            rom[21688] = 8'hcd ;
            rom[21689] = 8'h1e ;
            rom[21690] = 8'h0e ;
            rom[21691] = 8'hd5 ;
            rom[21692] = 8'he5 ;
            rom[21693] = 8'hde ;
            rom[21694] = 8'h1f ;
            rom[21695] = 8'hd7 ;
            rom[21696] = 8'ha2 ;
            rom[21697] = 8'h15 ;
            rom[21698] = 8'hf3 ;
            rom[21699] = 8'h18 ;
            rom[21700] = 8'h25 ;
            rom[21701] = 8'h05 ;
            rom[21702] = 8'hf8 ;
            rom[21703] = 8'he0 ;
            rom[21704] = 8'h0a ;
            rom[21705] = 8'h00 ;
            rom[21706] = 8'h0f ;
            rom[21707] = 8'h14 ;
            rom[21708] = 8'h08 ;
            rom[21709] = 8'heb ;
            rom[21710] = 8'h17 ;
            rom[21711] = 8'h11 ;
            rom[21712] = 8'hfa ;
            rom[21713] = 8'hbb ;
            rom[21714] = 8'hfa ;
            rom[21715] = 8'h04 ;
            rom[21716] = 8'hd2 ;
            rom[21717] = 8'hfd ;
            rom[21718] = 8'he8 ;
            rom[21719] = 8'h19 ;
            rom[21720] = 8'h01 ;
            rom[21721] = 8'hf0 ;
            rom[21722] = 8'h29 ;
            rom[21723] = 8'h11 ;
            rom[21724] = 8'h1c ;
            rom[21725] = 8'h16 ;
            rom[21726] = 8'h1b ;
            rom[21727] = 8'h06 ;
            rom[21728] = 8'heb ;
            rom[21729] = 8'he2 ;
            rom[21730] = 8'hfe ;
            rom[21731] = 8'hfb ;
            rom[21732] = 8'hb3 ;
            rom[21733] = 8'h04 ;
            rom[21734] = 8'hf7 ;
            rom[21735] = 8'he6 ;
            rom[21736] = 8'hd1 ;
            rom[21737] = 8'hd0 ;
            rom[21738] = 8'h02 ;
            rom[21739] = 8'h11 ;
            rom[21740] = 8'h27 ;
            rom[21741] = 8'h07 ;
            rom[21742] = 8'h21 ;
            rom[21743] = 8'he1 ;
            rom[21744] = 8'he8 ;
            rom[21745] = 8'hf0 ;
            rom[21746] = 8'h1c ;
            rom[21747] = 8'hd7 ;
            rom[21748] = 8'h17 ;
            rom[21749] = 8'h03 ;
            rom[21750] = 8'hf6 ;
            rom[21751] = 8'h01 ;
            rom[21752] = 8'hf6 ;
            rom[21753] = 8'hc0 ;
            rom[21754] = 8'hf0 ;
            rom[21755] = 8'he8 ;
            rom[21756] = 8'he0 ;
            rom[21757] = 8'hd8 ;
            rom[21758] = 8'hd9 ;
            rom[21759] = 8'hf1 ;
            rom[21760] = 8'hd9 ;
            rom[21761] = 8'h14 ;
            rom[21762] = 8'hf6 ;
            rom[21763] = 8'h07 ;
            rom[21764] = 8'h09 ;
            rom[21765] = 8'h02 ;
            rom[21766] = 8'h01 ;
            rom[21767] = 8'hf0 ;
            rom[21768] = 8'h0b ;
            rom[21769] = 8'hd8 ;
            rom[21770] = 8'h08 ;
            rom[21771] = 8'hf2 ;
            rom[21772] = 8'hf1 ;
            rom[21773] = 8'h12 ;
            rom[21774] = 8'h0e ;
            rom[21775] = 8'hf6 ;
            rom[21776] = 8'h14 ;
            rom[21777] = 8'h2d ;
            rom[21778] = 8'hcc ;
            rom[21779] = 8'hf4 ;
            rom[21780] = 8'h12 ;
            rom[21781] = 8'hfc ;
            rom[21782] = 8'hea ;
            rom[21783] = 8'hfd ;
            rom[21784] = 8'h04 ;
            rom[21785] = 8'hf1 ;
            rom[21786] = 8'h16 ;
            rom[21787] = 8'he6 ;
            rom[21788] = 8'hfc ;
            rom[21789] = 8'hc6 ;
            rom[21790] = 8'hd9 ;
            rom[21791] = 8'hc6 ;
            rom[21792] = 8'h1a ;
            rom[21793] = 8'hf7 ;
            rom[21794] = 8'hfa ;
            rom[21795] = 8'h10 ;
            rom[21796] = 8'hdf ;
            rom[21797] = 8'h10 ;
            rom[21798] = 8'he4 ;
            rom[21799] = 8'h0e ;
            rom[21800] = 8'hdc ;
            rom[21801] = 8'hee ;
            rom[21802] = 8'h07 ;
            rom[21803] = 8'h17 ;
            rom[21804] = 8'h18 ;
            rom[21805] = 8'h08 ;
            rom[21806] = 8'he9 ;
            rom[21807] = 8'hf2 ;
            rom[21808] = 8'hef ;
            rom[21809] = 8'hf1 ;
            rom[21810] = 8'hf9 ;
            rom[21811] = 8'hce ;
            rom[21812] = 8'hf8 ;
            rom[21813] = 8'hff ;
            rom[21814] = 8'hf8 ;
            rom[21815] = 8'h06 ;
            rom[21816] = 8'h03 ;
            rom[21817] = 8'hf0 ;
            rom[21818] = 8'hf4 ;
            rom[21819] = 8'hed ;
            rom[21820] = 8'h0e ;
            rom[21821] = 8'h03 ;
            rom[21822] = 8'h17 ;
            rom[21823] = 8'hfc ;
            rom[21824] = 8'he7 ;
            rom[21825] = 8'hb5 ;
            rom[21826] = 8'hf8 ;
            rom[21827] = 8'hf6 ;
            rom[21828] = 8'hef ;
            rom[21829] = 8'h07 ;
            rom[21830] = 8'hea ;
            rom[21831] = 8'h08 ;
            rom[21832] = 8'h05 ;
            rom[21833] = 8'hf7 ;
            rom[21834] = 8'hf1 ;
            rom[21835] = 8'hf4 ;
            rom[21836] = 8'h11 ;
            rom[21837] = 8'hd4 ;
            rom[21838] = 8'hf4 ;
            rom[21839] = 8'he7 ;
            rom[21840] = 8'h1e ;
            rom[21841] = 8'hfe ;
            rom[21842] = 8'hf2 ;
            rom[21843] = 8'h08 ;
            rom[21844] = 8'hec ;
            rom[21845] = 8'hde ;
            rom[21846] = 8'h05 ;
            rom[21847] = 8'he9 ;
            rom[21848] = 8'he6 ;
            rom[21849] = 8'hf3 ;
            rom[21850] = 8'hf8 ;
            rom[21851] = 8'h06 ;
            rom[21852] = 8'h13 ;
            rom[21853] = 8'h0f ;
            rom[21854] = 8'hf5 ;
            rom[21855] = 8'h09 ;
            rom[21856] = 8'hc3 ;
            rom[21857] = 8'h07 ;
            rom[21858] = 8'h02 ;
            rom[21859] = 8'h1c ;
            rom[21860] = 8'hfa ;
            rom[21861] = 8'hf5 ;
            rom[21862] = 8'h20 ;
            rom[21863] = 8'he4 ;
            rom[21864] = 8'h1a ;
            rom[21865] = 8'h20 ;
            rom[21866] = 8'h0d ;
            rom[21867] = 8'hfa ;
            rom[21868] = 8'hff ;
            rom[21869] = 8'hfc ;
            rom[21870] = 8'hcb ;
            rom[21871] = 8'hf4 ;
            rom[21872] = 8'h24 ;
            rom[21873] = 8'h1c ;
            rom[21874] = 8'h28 ;
            rom[21875] = 8'hf6 ;
            rom[21876] = 8'h02 ;
            rom[21877] = 8'hda ;
            rom[21878] = 8'h0f ;
            rom[21879] = 8'h19 ;
            rom[21880] = 8'hc5 ;
            rom[21881] = 8'h05 ;
            rom[21882] = 8'h0f ;
            rom[21883] = 8'hee ;
            rom[21884] = 8'he6 ;
            rom[21885] = 8'h11 ;
            rom[21886] = 8'h0d ;
            rom[21887] = 8'h04 ;
            rom[21888] = 8'h10 ;
            rom[21889] = 8'hf2 ;
            rom[21890] = 8'hfc ;
            rom[21891] = 8'h08 ;
            rom[21892] = 8'h18 ;
            rom[21893] = 8'hf2 ;
            rom[21894] = 8'h0c ;
            rom[21895] = 8'hd9 ;
            rom[21896] = 8'hd9 ;
            rom[21897] = 8'hdf ;
            rom[21898] = 8'h32 ;
            rom[21899] = 8'h05 ;
            rom[21900] = 8'h0c ;
            rom[21901] = 8'hf5 ;
            rom[21902] = 8'hc1 ;
            rom[21903] = 8'h00 ;
            rom[21904] = 8'hd9 ;
            rom[21905] = 8'hf7 ;
            rom[21906] = 8'hf9 ;
            rom[21907] = 8'he8 ;
            rom[21908] = 8'hef ;
            rom[21909] = 8'hf6 ;
            rom[21910] = 8'h0f ;
            rom[21911] = 8'hc1 ;
            rom[21912] = 8'h01 ;
            rom[21913] = 8'heb ;
            rom[21914] = 8'he5 ;
            rom[21915] = 8'he9 ;
            rom[21916] = 8'hfd ;
            rom[21917] = 8'hd7 ;
            rom[21918] = 8'h08 ;
            rom[21919] = 8'hfd ;
            rom[21920] = 8'h19 ;
            rom[21921] = 8'h18 ;
            rom[21922] = 8'hf8 ;
            rom[21923] = 8'h14 ;
            rom[21924] = 8'he9 ;
            rom[21925] = 8'h00 ;
            rom[21926] = 8'hc6 ;
            rom[21927] = 8'h11 ;
            rom[21928] = 8'hfc ;
            rom[21929] = 8'hf9 ;
            rom[21930] = 8'h0b ;
            rom[21931] = 8'hf8 ;
            rom[21932] = 8'h14 ;
            rom[21933] = 8'h03 ;
            rom[21934] = 8'hf7 ;
            rom[21935] = 8'h03 ;
            rom[21936] = 8'h14 ;
            rom[21937] = 8'hea ;
            rom[21938] = 8'hfe ;
            rom[21939] = 8'h05 ;
            rom[21940] = 8'h08 ;
            rom[21941] = 8'h00 ;
            rom[21942] = 8'hed ;
            rom[21943] = 8'h1d ;
            rom[21944] = 8'h0c ;
            rom[21945] = 8'hfe ;
            rom[21946] = 8'hf6 ;
            rom[21947] = 8'he4 ;
            rom[21948] = 8'hf6 ;
            rom[21949] = 8'hfb ;
            rom[21950] = 8'hde ;
            rom[21951] = 8'hd5 ;
            rom[21952] = 8'hf2 ;
            rom[21953] = 8'hdf ;
            rom[21954] = 8'hf4 ;
            rom[21955] = 8'h1d ;
            rom[21956] = 8'hdb ;
            rom[21957] = 8'he1 ;
            rom[21958] = 8'hec ;
            rom[21959] = 8'h03 ;
            rom[21960] = 8'h06 ;
            rom[21961] = 8'he4 ;
            rom[21962] = 8'hff ;
            rom[21963] = 8'h0c ;
            rom[21964] = 8'hfa ;
            rom[21965] = 8'hed ;
            rom[21966] = 8'hf0 ;
            rom[21967] = 8'he8 ;
            rom[21968] = 8'hfb ;
            rom[21969] = 8'hf1 ;
            rom[21970] = 8'he4 ;
            rom[21971] = 8'hfe ;
            rom[21972] = 8'hf4 ;
            rom[21973] = 8'hde ;
            rom[21974] = 8'h03 ;
            rom[21975] = 8'h18 ;
            rom[21976] = 8'he6 ;
            rom[21977] = 8'h0a ;
            rom[21978] = 8'h1f ;
            rom[21979] = 8'h29 ;
            rom[21980] = 8'h10 ;
            rom[21981] = 8'hc7 ;
            rom[21982] = 8'h1f ;
            rom[21983] = 8'hdb ;
            rom[21984] = 8'hee ;
            rom[21985] = 8'h09 ;
            rom[21986] = 8'hfd ;
            rom[21987] = 8'hf1 ;
            rom[21988] = 8'hfb ;
            rom[21989] = 8'hee ;
            rom[21990] = 8'h06 ;
            rom[21991] = 8'he8 ;
            rom[21992] = 8'hfe ;
            rom[21993] = 8'h13 ;
            rom[21994] = 8'hcd ;
            rom[21995] = 8'hf1 ;
            rom[21996] = 8'h00 ;
            rom[21997] = 8'h0d ;
            rom[21998] = 8'hee ;
            rom[21999] = 8'h08 ;
            rom[22000] = 8'hdd ;
            rom[22001] = 8'h15 ;
            rom[22002] = 8'h1a ;
            rom[22003] = 8'hf9 ;
            rom[22004] = 8'he1 ;
            rom[22005] = 8'h0b ;
            rom[22006] = 8'h01 ;
            rom[22007] = 8'hef ;
            rom[22008] = 8'hfe ;
            rom[22009] = 8'hd8 ;
            rom[22010] = 8'h1e ;
            rom[22011] = 8'h04 ;
            rom[22012] = 8'hfd ;
            rom[22013] = 8'hfc ;
            rom[22014] = 8'h06 ;
            rom[22015] = 8'hf8 ;
            rom[22016] = 8'h12 ;
            rom[22017] = 8'he0 ;
            rom[22018] = 8'h0b ;
            rom[22019] = 8'h1b ;
            rom[22020] = 8'hde ;
            rom[22021] = 8'hf9 ;
            rom[22022] = 8'hc5 ;
            rom[22023] = 8'hf3 ;
            rom[22024] = 8'hef ;
            rom[22025] = 8'h06 ;
            rom[22026] = 8'he6 ;
            rom[22027] = 8'h10 ;
            rom[22028] = 8'hef ;
            rom[22029] = 8'h19 ;
            rom[22030] = 8'h03 ;
            rom[22031] = 8'hf7 ;
            rom[22032] = 8'h20 ;
            rom[22033] = 8'h0e ;
            rom[22034] = 8'hcd ;
            rom[22035] = 8'h1c ;
            rom[22036] = 8'h0a ;
            rom[22037] = 8'he5 ;
            rom[22038] = 8'hed ;
            rom[22039] = 8'hdd ;
            rom[22040] = 8'hf4 ;
            rom[22041] = 8'hfd ;
            rom[22042] = 8'h09 ;
            rom[22043] = 8'hb6 ;
            rom[22044] = 8'he9 ;
            rom[22045] = 8'hee ;
            rom[22046] = 8'h02 ;
            rom[22047] = 8'h1e ;
            rom[22048] = 8'hf7 ;
            rom[22049] = 8'h0d ;
            rom[22050] = 8'h05 ;
            rom[22051] = 8'hf5 ;
            rom[22052] = 8'hbf ;
            rom[22053] = 8'hf0 ;
            rom[22054] = 8'hfe ;
            rom[22055] = 8'hda ;
            rom[22056] = 8'he2 ;
            rom[22057] = 8'hc0 ;
            rom[22058] = 8'h0d ;
            rom[22059] = 8'hfd ;
            rom[22060] = 8'h18 ;
            rom[22061] = 8'h03 ;
            rom[22062] = 8'hd4 ;
            rom[22063] = 8'h10 ;
            rom[22064] = 8'hd8 ;
            rom[22065] = 8'hf0 ;
            rom[22066] = 8'h0c ;
            rom[22067] = 8'hf8 ;
            rom[22068] = 8'hf8 ;
            rom[22069] = 8'hfe ;
            rom[22070] = 8'hff ;
            rom[22071] = 8'hf1 ;
            rom[22072] = 8'h13 ;
            rom[22073] = 8'hcd ;
            rom[22074] = 8'h09 ;
            rom[22075] = 8'hdc ;
            rom[22076] = 8'hce ;
            rom[22077] = 8'he3 ;
            rom[22078] = 8'h08 ;
            rom[22079] = 8'hdf ;
            rom[22080] = 8'hed ;
            rom[22081] = 8'h0a ;
            rom[22082] = 8'hfb ;
            rom[22083] = 8'hbc ;
            rom[22084] = 8'he9 ;
            rom[22085] = 8'hdb ;
            rom[22086] = 8'hd3 ;
            rom[22087] = 8'h0d ;
            rom[22088] = 8'h07 ;
            rom[22089] = 8'h07 ;
            rom[22090] = 8'he4 ;
            rom[22091] = 8'hdc ;
            rom[22092] = 8'hf8 ;
            rom[22093] = 8'h00 ;
            rom[22094] = 8'h02 ;
            rom[22095] = 8'hfe ;
            rom[22096] = 8'hf4 ;
            rom[22097] = 8'h0f ;
            rom[22098] = 8'h07 ;
            rom[22099] = 8'hf4 ;
            rom[22100] = 8'hf1 ;
            rom[22101] = 8'h0a ;
            rom[22102] = 8'h1a ;
            rom[22103] = 8'he0 ;
            rom[22104] = 8'h05 ;
            rom[22105] = 8'hf3 ;
            rom[22106] = 8'h24 ;
            rom[22107] = 8'h15 ;
            rom[22108] = 8'hf1 ;
            rom[22109] = 8'hec ;
            rom[22110] = 8'h06 ;
            rom[22111] = 8'he4 ;
            rom[22112] = 8'h12 ;
            rom[22113] = 8'he7 ;
            rom[22114] = 8'h13 ;
            rom[22115] = 8'h0c ;
            rom[22116] = 8'hca ;
            rom[22117] = 8'heb ;
            rom[22118] = 8'h07 ;
            rom[22119] = 8'h16 ;
            rom[22120] = 8'h01 ;
            rom[22121] = 8'h0d ;
            rom[22122] = 8'he2 ;
            rom[22123] = 8'hfd ;
            rom[22124] = 8'h09 ;
            rom[22125] = 8'h15 ;
            rom[22126] = 8'h04 ;
            rom[22127] = 8'h0e ;
            rom[22128] = 8'he9 ;
            rom[22129] = 8'he7 ;
            rom[22130] = 8'hfb ;
            rom[22131] = 8'hfc ;
            rom[22132] = 8'hef ;
            rom[22133] = 8'he6 ;
            rom[22134] = 8'hef ;
            rom[22135] = 8'h01 ;
            rom[22136] = 8'h0a ;
            rom[22137] = 8'h05 ;
            rom[22138] = 8'he7 ;
            rom[22139] = 8'he2 ;
            rom[22140] = 8'hce ;
            rom[22141] = 8'he6 ;
            rom[22142] = 8'h00 ;
            rom[22143] = 8'h2c ;
            rom[22144] = 8'h04 ;
            rom[22145] = 8'he9 ;
            rom[22146] = 8'h01 ;
            rom[22147] = 8'hfb ;
            rom[22148] = 8'h0d ;
            rom[22149] = 8'h01 ;
            rom[22150] = 8'h01 ;
            rom[22151] = 8'he4 ;
            rom[22152] = 8'hcb ;
            rom[22153] = 8'h00 ;
            rom[22154] = 8'hec ;
            rom[22155] = 8'h0d ;
            rom[22156] = 8'he7 ;
            rom[22157] = 8'h0b ;
            rom[22158] = 8'hd0 ;
            rom[22159] = 8'hca ;
            rom[22160] = 8'h0c ;
            rom[22161] = 8'h09 ;
            rom[22162] = 8'he0 ;
            rom[22163] = 8'hfc ;
            rom[22164] = 8'h10 ;
            rom[22165] = 8'hed ;
            rom[22166] = 8'h03 ;
            rom[22167] = 8'h90 ;
            rom[22168] = 8'he8 ;
            rom[22169] = 8'h0f ;
            rom[22170] = 8'hf1 ;
            rom[22171] = 8'hd0 ;
            rom[22172] = 8'he7 ;
            rom[22173] = 8'hd5 ;
            rom[22174] = 8'hee ;
            rom[22175] = 8'h1a ;
            rom[22176] = 8'hf6 ;
            rom[22177] = 8'h2f ;
            rom[22178] = 8'h00 ;
            rom[22179] = 8'hdd ;
            rom[22180] = 8'h15 ;
            rom[22181] = 8'hfd ;
            rom[22182] = 8'he4 ;
            rom[22183] = 8'h1f ;
            rom[22184] = 8'hf3 ;
            rom[22185] = 8'hf4 ;
            rom[22186] = 8'h14 ;
            rom[22187] = 8'hec ;
            rom[22188] = 8'hee ;
            rom[22189] = 8'h10 ;
            rom[22190] = 8'hd8 ;
            rom[22191] = 8'hf3 ;
            rom[22192] = 8'h16 ;
            rom[22193] = 8'he8 ;
            rom[22194] = 8'he9 ;
            rom[22195] = 8'h01 ;
            rom[22196] = 8'h16 ;
            rom[22197] = 8'hea ;
            rom[22198] = 8'hef ;
            rom[22199] = 8'he9 ;
            rom[22200] = 8'he9 ;
            rom[22201] = 8'he4 ;
            rom[22202] = 8'hdb ;
            rom[22203] = 8'h11 ;
            rom[22204] = 8'hfe ;
            rom[22205] = 8'h0c ;
            rom[22206] = 8'h0f ;
            rom[22207] = 8'hda ;
            rom[22208] = 8'h05 ;
            rom[22209] = 8'hff ;
            rom[22210] = 8'h0c ;
            rom[22211] = 8'hd4 ;
            rom[22212] = 8'hed ;
            rom[22213] = 8'h0f ;
            rom[22214] = 8'hf4 ;
            rom[22215] = 8'h19 ;
            rom[22216] = 8'hf4 ;
            rom[22217] = 8'hec ;
            rom[22218] = 8'hff ;
            rom[22219] = 8'hde ;
            rom[22220] = 8'h11 ;
            rom[22221] = 8'h16 ;
            rom[22222] = 8'hed ;
            rom[22223] = 8'hf8 ;
            rom[22224] = 8'hdd ;
            rom[22225] = 8'hde ;
            rom[22226] = 8'h00 ;
            rom[22227] = 8'hf4 ;
            rom[22228] = 8'hd4 ;
            rom[22229] = 8'hdc ;
            rom[22230] = 8'h05 ;
            rom[22231] = 8'h23 ;
            rom[22232] = 8'hfb ;
            rom[22233] = 8'hec ;
            rom[22234] = 8'h14 ;
            rom[22235] = 8'h0e ;
            rom[22236] = 8'hc2 ;
            rom[22237] = 8'hd2 ;
            rom[22238] = 8'h1a ;
            rom[22239] = 8'h07 ;
            rom[22240] = 8'hf6 ;
            rom[22241] = 8'hfe ;
            rom[22242] = 8'hff ;
            rom[22243] = 8'hf3 ;
            rom[22244] = 8'hea ;
            rom[22245] = 8'h0b ;
            rom[22246] = 8'h18 ;
            rom[22247] = 8'hff ;
            rom[22248] = 8'hde ;
            rom[22249] = 8'h03 ;
            rom[22250] = 8'hd5 ;
            rom[22251] = 8'hc7 ;
            rom[22252] = 8'h1d ;
            rom[22253] = 8'h03 ;
            rom[22254] = 8'h00 ;
            rom[22255] = 8'h1a ;
            rom[22256] = 8'h04 ;
            rom[22257] = 8'h0d ;
            rom[22258] = 8'h10 ;
            rom[22259] = 8'hd2 ;
            rom[22260] = 8'heb ;
            rom[22261] = 8'h0d ;
            rom[22262] = 8'hf8 ;
            rom[22263] = 8'h11 ;
            rom[22264] = 8'h1a ;
            rom[22265] = 8'h06 ;
            rom[22266] = 8'h11 ;
            rom[22267] = 8'hf8 ;
            rom[22268] = 8'hcd ;
            rom[22269] = 8'hfd ;
            rom[22270] = 8'h01 ;
            rom[22271] = 8'h0b ;
            rom[22272] = 8'hea ;
            rom[22273] = 8'h05 ;
            rom[22274] = 8'h02 ;
            rom[22275] = 8'he4 ;
            rom[22276] = 8'he7 ;
            rom[22277] = 8'hdb ;
            rom[22278] = 8'hff ;
            rom[22279] = 8'h06 ;
            rom[22280] = 8'he6 ;
            rom[22281] = 8'h14 ;
            rom[22282] = 8'h16 ;
            rom[22283] = 8'h0f ;
            rom[22284] = 8'hef ;
            rom[22285] = 8'h10 ;
            rom[22286] = 8'hfb ;
            rom[22287] = 8'he4 ;
            rom[22288] = 8'hd4 ;
            rom[22289] = 8'hf9 ;
            rom[22290] = 8'h12 ;
            rom[22291] = 8'hea ;
            rom[22292] = 8'he9 ;
            rom[22293] = 8'hec ;
            rom[22294] = 8'hf1 ;
            rom[22295] = 8'h03 ;
            rom[22296] = 8'he7 ;
            rom[22297] = 8'h08 ;
            rom[22298] = 8'hee ;
            rom[22299] = 8'hf8 ;
            rom[22300] = 8'hf8 ;
            rom[22301] = 8'h18 ;
            rom[22302] = 8'h15 ;
            rom[22303] = 8'h03 ;
            rom[22304] = 8'hb8 ;
            rom[22305] = 8'hd5 ;
            rom[22306] = 8'hf8 ;
            rom[22307] = 8'h06 ;
            rom[22308] = 8'h1b ;
            rom[22309] = 8'hc8 ;
            rom[22310] = 8'h13 ;
            rom[22311] = 8'hf7 ;
            rom[22312] = 8'h2b ;
            rom[22313] = 8'hf7 ;
            rom[22314] = 8'hf5 ;
            rom[22315] = 8'hce ;
            rom[22316] = 8'hc7 ;
            rom[22317] = 8'hc9 ;
            rom[22318] = 8'h25 ;
            rom[22319] = 8'hf3 ;
            rom[22320] = 8'h01 ;
            rom[22321] = 8'hd0 ;
            rom[22322] = 8'he9 ;
            rom[22323] = 8'h24 ;
            rom[22324] = 8'hf3 ;
            rom[22325] = 8'hf3 ;
            rom[22326] = 8'hf8 ;
            rom[22327] = 8'h0a ;
            rom[22328] = 8'hcd ;
            rom[22329] = 8'h0f ;
            rom[22330] = 8'h33 ;
            rom[22331] = 8'h03 ;
            rom[22332] = 8'hfb ;
            rom[22333] = 8'hfb ;
            rom[22334] = 8'hdb ;
            rom[22335] = 8'h25 ;
            rom[22336] = 8'hf6 ;
            rom[22337] = 8'hf7 ;
            rom[22338] = 8'hfe ;
            rom[22339] = 8'he4 ;
            rom[22340] = 8'h1d ;
            rom[22341] = 8'h03 ;
            rom[22342] = 8'h05 ;
            rom[22343] = 8'hf7 ;
            rom[22344] = 8'h04 ;
            rom[22345] = 8'h0f ;
            rom[22346] = 8'h00 ;
            rom[22347] = 8'h1b ;
            rom[22348] = 8'hb7 ;
            rom[22349] = 8'h02 ;
            rom[22350] = 8'hfc ;
            rom[22351] = 8'hf9 ;
            rom[22352] = 8'hf7 ;
            rom[22353] = 8'hf5 ;
            rom[22354] = 8'hc5 ;
            rom[22355] = 8'he0 ;
            rom[22356] = 8'h09 ;
            rom[22357] = 8'h07 ;
            rom[22358] = 8'hc8 ;
            rom[22359] = 8'h12 ;
            rom[22360] = 8'h10 ;
            rom[22361] = 8'he4 ;
            rom[22362] = 8'hd9 ;
            rom[22363] = 8'hce ;
            rom[22364] = 8'hea ;
            rom[22365] = 8'he6 ;
            rom[22366] = 8'hef ;
            rom[22367] = 8'h1c ;
            rom[22368] = 8'h24 ;
            rom[22369] = 8'hf0 ;
            rom[22370] = 8'hf1 ;
            rom[22371] = 8'hec ;
            rom[22372] = 8'h1e ;
            rom[22373] = 8'hdd ;
            rom[22374] = 8'hff ;
            rom[22375] = 8'h0e ;
            rom[22376] = 8'he6 ;
            rom[22377] = 8'hd9 ;
            rom[22378] = 8'he1 ;
            rom[22379] = 8'h21 ;
            rom[22380] = 8'hf8 ;
            rom[22381] = 8'he6 ;
            rom[22382] = 8'h0f ;
            rom[22383] = 8'hfd ;
            rom[22384] = 8'h0d ;
            rom[22385] = 8'hfb ;
            rom[22386] = 8'hf3 ;
            rom[22387] = 8'hf6 ;
            rom[22388] = 8'h00 ;
            rom[22389] = 8'hfd ;
            rom[22390] = 8'h2c ;
            rom[22391] = 8'hce ;
            rom[22392] = 8'hdb ;
            rom[22393] = 8'h11 ;
            rom[22394] = 8'h11 ;
            rom[22395] = 8'h13 ;
            rom[22396] = 8'h12 ;
            rom[22397] = 8'hbe ;
            rom[22398] = 8'heb ;
            rom[22399] = 8'he0 ;
            rom[22400] = 8'hd6 ;
            rom[22401] = 8'h0c ;
            rom[22402] = 8'hf7 ;
            rom[22403] = 8'hec ;
            rom[22404] = 8'hea ;
            rom[22405] = 8'hed ;
            rom[22406] = 8'h08 ;
            rom[22407] = 8'h1b ;
            rom[22408] = 8'h10 ;
            rom[22409] = 8'h00 ;
            rom[22410] = 8'hc8 ;
            rom[22411] = 8'hfd ;
            rom[22412] = 8'hfc ;
            rom[22413] = 8'h17 ;
            rom[22414] = 8'h09 ;
            rom[22415] = 8'h19 ;
            rom[22416] = 8'h27 ;
            rom[22417] = 8'h1a ;
            rom[22418] = 8'hfd ;
            rom[22419] = 8'hf6 ;
            rom[22420] = 8'hf0 ;
            rom[22421] = 8'h06 ;
            rom[22422] = 8'h1e ;
            rom[22423] = 8'h25 ;
            rom[22424] = 8'h2d ;
            rom[22425] = 8'hfc ;
            rom[22426] = 8'h0b ;
            rom[22427] = 8'h0a ;
            rom[22428] = 8'hf0 ;
            rom[22429] = 8'h0f ;
            rom[22430] = 8'h07 ;
            rom[22431] = 8'h07 ;
            rom[22432] = 8'h1b ;
            rom[22433] = 8'h12 ;
            rom[22434] = 8'hf1 ;
            rom[22435] = 8'he7 ;
            rom[22436] = 8'hcb ;
            rom[22437] = 8'h01 ;
            rom[22438] = 8'h10 ;
            rom[22439] = 8'hde ;
            rom[22440] = 8'hdd ;
            rom[22441] = 8'hf3 ;
            rom[22442] = 8'hf0 ;
            rom[22443] = 8'h17 ;
            rom[22444] = 8'h24 ;
            rom[22445] = 8'hf1 ;
            rom[22446] = 8'hb5 ;
            rom[22447] = 8'hf1 ;
            rom[22448] = 8'he7 ;
            rom[22449] = 8'hfb ;
            rom[22450] = 8'h16 ;
            rom[22451] = 8'he7 ;
            rom[22452] = 8'hfd ;
            rom[22453] = 8'hdb ;
            rom[22454] = 8'hff ;
            rom[22455] = 8'h07 ;
            rom[22456] = 8'h0f ;
            rom[22457] = 8'h05 ;
            rom[22458] = 8'he2 ;
            rom[22459] = 8'hca ;
            rom[22460] = 8'h0c ;
            rom[22461] = 8'hf8 ;
            rom[22462] = 8'h17 ;
            rom[22463] = 8'h13 ;
            rom[22464] = 8'h1e ;
            rom[22465] = 8'hda ;
            rom[22466] = 8'he5 ;
            rom[22467] = 8'h21 ;
            rom[22468] = 8'h09 ;
            rom[22469] = 8'hf0 ;
            rom[22470] = 8'hf7 ;
            rom[22471] = 8'h01 ;
            rom[22472] = 8'hdc ;
            rom[22473] = 8'hf4 ;
            rom[22474] = 8'hd8 ;
            rom[22475] = 8'he0 ;
            rom[22476] = 8'h2a ;
            rom[22477] = 8'h16 ;
            rom[22478] = 8'hf0 ;
            rom[22479] = 8'h0e ;
            rom[22480] = 8'hf4 ;
            rom[22481] = 8'h23 ;
            rom[22482] = 8'h38 ;
            rom[22483] = 8'h1b ;
            rom[22484] = 8'h1c ;
            rom[22485] = 8'hee ;
            rom[22486] = 8'hdc ;
            rom[22487] = 8'hd4 ;
            rom[22488] = 8'hf9 ;
            rom[22489] = 8'h1a ;
            rom[22490] = 8'he0 ;
            rom[22491] = 8'hf6 ;
            rom[22492] = 8'h01 ;
            rom[22493] = 8'h27 ;
            rom[22494] = 8'hf4 ;
            rom[22495] = 8'hff ;
            rom[22496] = 8'hfd ;
            rom[22497] = 8'h1c ;
            rom[22498] = 8'hc8 ;
            rom[22499] = 8'h33 ;
            rom[22500] = 8'h18 ;
            rom[22501] = 8'h13 ;
            rom[22502] = 8'h0c ;
            rom[22503] = 8'hfb ;
            rom[22504] = 8'h34 ;
            rom[22505] = 8'hea ;
            rom[22506] = 8'hcc ;
            rom[22507] = 8'h0d ;
            rom[22508] = 8'he3 ;
            rom[22509] = 8'h1b ;
            rom[22510] = 8'he7 ;
            rom[22511] = 8'hdf ;
            rom[22512] = 8'h0e ;
            rom[22513] = 8'hf1 ;
            rom[22514] = 8'hb7 ;
            rom[22515] = 8'h15 ;
            rom[22516] = 8'hfc ;
            rom[22517] = 8'hec ;
            rom[22518] = 8'heb ;
            rom[22519] = 8'he8 ;
            rom[22520] = 8'hd9 ;
            rom[22521] = 8'h05 ;
            rom[22522] = 8'h00 ;
            rom[22523] = 8'h2a ;
            rom[22524] = 8'hfd ;
            rom[22525] = 8'h12 ;
            rom[22526] = 8'h0d ;
            rom[22527] = 8'h36 ;
            rom[22528] = 8'hd7 ;
            rom[22529] = 8'he5 ;
            rom[22530] = 8'he7 ;
            rom[22531] = 8'hf3 ;
            rom[22532] = 8'he1 ;
            rom[22533] = 8'h1a ;
            rom[22534] = 8'h0b ;
            rom[22535] = 8'hfd ;
            rom[22536] = 8'h18 ;
            rom[22537] = 8'h02 ;
            rom[22538] = 8'hee ;
            rom[22539] = 8'he7 ;
            rom[22540] = 8'hd6 ;
            rom[22541] = 8'hf0 ;
            rom[22542] = 8'h09 ;
            rom[22543] = 8'h0f ;
            rom[22544] = 8'h0d ;
            rom[22545] = 8'hda ;
            rom[22546] = 8'hc7 ;
            rom[22547] = 8'h0c ;
            rom[22548] = 8'hdf ;
            rom[22549] = 8'h1b ;
            rom[22550] = 8'h0b ;
            rom[22551] = 8'h05 ;
            rom[22552] = 8'hf7 ;
            rom[22553] = 8'h09 ;
            rom[22554] = 8'h07 ;
            rom[22555] = 8'h07 ;
            rom[22556] = 8'he8 ;
            rom[22557] = 8'hc8 ;
            rom[22558] = 8'he0 ;
            rom[22559] = 8'hfc ;
            rom[22560] = 8'hd9 ;
            rom[22561] = 8'hdf ;
            rom[22562] = 8'h05 ;
            rom[22563] = 8'h11 ;
            rom[22564] = 8'heb ;
            rom[22565] = 8'hec ;
            rom[22566] = 8'hae ;
            rom[22567] = 8'hf3 ;
            rom[22568] = 8'h02 ;
            rom[22569] = 8'hf8 ;
            rom[22570] = 8'hf7 ;
            rom[22571] = 8'h0b ;
            rom[22572] = 8'hf9 ;
            rom[22573] = 8'hff ;
            rom[22574] = 8'hbc ;
            rom[22575] = 8'hf1 ;
            rom[22576] = 8'hf1 ;
            rom[22577] = 8'h12 ;
            rom[22578] = 8'h13 ;
            rom[22579] = 8'haf ;
            rom[22580] = 8'h1a ;
            rom[22581] = 8'he1 ;
            rom[22582] = 8'hf5 ;
            rom[22583] = 8'h1c ;
            rom[22584] = 8'h16 ;
            rom[22585] = 8'he7 ;
            rom[22586] = 8'h05 ;
            rom[22587] = 8'he7 ;
            rom[22588] = 8'hf3 ;
            rom[22589] = 8'hc7 ;
            rom[22590] = 8'h05 ;
            rom[22591] = 8'heb ;
            rom[22592] = 8'hf8 ;
            rom[22593] = 8'hee ;
            rom[22594] = 8'he3 ;
            rom[22595] = 8'h26 ;
            rom[22596] = 8'h03 ;
            rom[22597] = 8'hd0 ;
            rom[22598] = 8'h06 ;
            rom[22599] = 8'hf8 ;
            rom[22600] = 8'h01 ;
            rom[22601] = 8'hd6 ;
            rom[22602] = 8'hff ;
            rom[22603] = 8'h19 ;
            rom[22604] = 8'h15 ;
            rom[22605] = 8'h03 ;
            rom[22606] = 8'hef ;
            rom[22607] = 8'he4 ;
            rom[22608] = 8'hdf ;
            rom[22609] = 8'h18 ;
            rom[22610] = 8'hfe ;
            rom[22611] = 8'hf5 ;
            rom[22612] = 8'h0c ;
            rom[22613] = 8'h06 ;
            rom[22614] = 8'hdf ;
            rom[22615] = 8'hf0 ;
            rom[22616] = 8'hed ;
            rom[22617] = 8'hd9 ;
            rom[22618] = 8'h1a ;
            rom[22619] = 8'h1c ;
            rom[22620] = 8'hfd ;
            rom[22621] = 8'hce ;
            rom[22622] = 8'hf1 ;
            rom[22623] = 8'h0e ;
            rom[22624] = 8'hf6 ;
            rom[22625] = 8'h14 ;
            rom[22626] = 8'h0c ;
            rom[22627] = 8'h0e ;
            rom[22628] = 8'hfc ;
            rom[22629] = 8'hce ;
            rom[22630] = 8'h1a ;
            rom[22631] = 8'hf8 ;
            rom[22632] = 8'h14 ;
            rom[22633] = 8'h15 ;
            rom[22634] = 8'hbc ;
            rom[22635] = 8'hf3 ;
            rom[22636] = 8'h04 ;
            rom[22637] = 8'h22 ;
            rom[22638] = 8'he5 ;
            rom[22639] = 8'hef ;
            rom[22640] = 8'hfb ;
            rom[22641] = 8'h03 ;
            rom[22642] = 8'hf5 ;
            rom[22643] = 8'hf8 ;
            rom[22644] = 8'he8 ;
            rom[22645] = 8'hd3 ;
            rom[22646] = 8'h01 ;
            rom[22647] = 8'h05 ;
            rom[22648] = 8'hf0 ;
            rom[22649] = 8'hff ;
            rom[22650] = 8'h1e ;
            rom[22651] = 8'h09 ;
            rom[22652] = 8'hdd ;
            rom[22653] = 8'he1 ;
            rom[22654] = 8'h03 ;
            rom[22655] = 8'hf1 ;
            rom[22656] = 8'he6 ;
            rom[22657] = 8'hdb ;
            rom[22658] = 8'h06 ;
            rom[22659] = 8'h1e ;
            rom[22660] = 8'hd1 ;
            rom[22661] = 8'h09 ;
            rom[22662] = 8'hcb ;
            rom[22663] = 8'h0f ;
            rom[22664] = 8'h16 ;
            rom[22665] = 8'h1e ;
            rom[22666] = 8'hf0 ;
            rom[22667] = 8'h38 ;
            rom[22668] = 8'h07 ;
            rom[22669] = 8'he3 ;
            rom[22670] = 8'h25 ;
            rom[22671] = 8'hef ;
            rom[22672] = 8'hf9 ;
            rom[22673] = 8'h0d ;
            rom[22674] = 8'hdc ;
            rom[22675] = 8'h01 ;
            rom[22676] = 8'h44 ;
            rom[22677] = 8'hf7 ;
            rom[22678] = 8'hfa ;
            rom[22679] = 8'h09 ;
            rom[22680] = 8'hfb ;
            rom[22681] = 8'h0e ;
            rom[22682] = 8'hfd ;
            rom[22683] = 8'hf4 ;
            rom[22684] = 8'hdf ;
            rom[22685] = 8'h0d ;
            rom[22686] = 8'h04 ;
            rom[22687] = 8'h04 ;
            rom[22688] = 8'heb ;
            rom[22689] = 8'hf0 ;
            rom[22690] = 8'hf7 ;
            rom[22691] = 8'he1 ;
            rom[22692] = 8'h0c ;
            rom[22693] = 8'h07 ;
            rom[22694] = 8'h06 ;
            rom[22695] = 8'hd6 ;
            rom[22696] = 8'h12 ;
            rom[22697] = 8'hc3 ;
            rom[22698] = 8'heb ;
            rom[22699] = 8'h02 ;
            rom[22700] = 8'hea ;
            rom[22701] = 8'hf5 ;
            rom[22702] = 8'hb2 ;
            rom[22703] = 8'he6 ;
            rom[22704] = 8'hce ;
            rom[22705] = 8'hfa ;
            rom[22706] = 8'h12 ;
            rom[22707] = 8'hf0 ;
            rom[22708] = 8'h01 ;
            rom[22709] = 8'hd4 ;
            rom[22710] = 8'h0a ;
            rom[22711] = 8'hf4 ;
            rom[22712] = 8'hfa ;
            rom[22713] = 8'hfd ;
            rom[22714] = 8'h1a ;
            rom[22715] = 8'hf6 ;
            rom[22716] = 8'h1b ;
            rom[22717] = 8'hce ;
            rom[22718] = 8'hef ;
            rom[22719] = 8'h00 ;
            rom[22720] = 8'hf4 ;
            rom[22721] = 8'hea ;
            rom[22722] = 8'h29 ;
            rom[22723] = 8'h09 ;
            rom[22724] = 8'h21 ;
            rom[22725] = 8'hfd ;
            rom[22726] = 8'hfb ;
            rom[22727] = 8'hfb ;
            rom[22728] = 8'he3 ;
            rom[22729] = 8'h16 ;
            rom[22730] = 8'h07 ;
            rom[22731] = 8'hfe ;
            rom[22732] = 8'h07 ;
            rom[22733] = 8'hea ;
            rom[22734] = 8'h15 ;
            rom[22735] = 8'hc7 ;
            rom[22736] = 8'he3 ;
            rom[22737] = 8'hf3 ;
            rom[22738] = 8'h19 ;
            rom[22739] = 8'hdb ;
            rom[22740] = 8'hf9 ;
            rom[22741] = 8'h0d ;
            rom[22742] = 8'hf9 ;
            rom[22743] = 8'hbb ;
            rom[22744] = 8'h33 ;
            rom[22745] = 8'he0 ;
            rom[22746] = 8'h23 ;
            rom[22747] = 8'h16 ;
            rom[22748] = 8'h19 ;
            rom[22749] = 8'hea ;
            rom[22750] = 8'hf5 ;
            rom[22751] = 8'hf7 ;
            rom[22752] = 8'hdf ;
            rom[22753] = 8'h16 ;
            rom[22754] = 8'hf9 ;
            rom[22755] = 8'h01 ;
            rom[22756] = 8'h04 ;
            rom[22757] = 8'h06 ;
            rom[22758] = 8'h1f ;
            rom[22759] = 8'h02 ;
            rom[22760] = 8'h04 ;
            rom[22761] = 8'h11 ;
            rom[22762] = 8'h13 ;
            rom[22763] = 8'hf0 ;
            rom[22764] = 8'h1c ;
            rom[22765] = 8'h03 ;
            rom[22766] = 8'hee ;
            rom[22767] = 8'hfb ;
            rom[22768] = 8'h03 ;
            rom[22769] = 8'hf8 ;
            rom[22770] = 8'h0f ;
            rom[22771] = 8'he1 ;
            rom[22772] = 8'h07 ;
            rom[22773] = 8'hdd ;
            rom[22774] = 8'h03 ;
            rom[22775] = 8'hfa ;
            rom[22776] = 8'he7 ;
            rom[22777] = 8'h24 ;
            rom[22778] = 8'h1e ;
            rom[22779] = 8'hf4 ;
            rom[22780] = 8'hcd ;
            rom[22781] = 8'h07 ;
            rom[22782] = 8'he4 ;
            rom[22783] = 8'h0e ;
            rom[22784] = 8'h03 ;
            rom[22785] = 8'hf8 ;
            rom[22786] = 8'h19 ;
            rom[22787] = 8'hf9 ;
            rom[22788] = 8'hf4 ;
            rom[22789] = 8'he9 ;
            rom[22790] = 8'h22 ;
            rom[22791] = 8'hed ;
            rom[22792] = 8'hf5 ;
            rom[22793] = 8'h02 ;
            rom[22794] = 8'h15 ;
            rom[22795] = 8'hf0 ;
            rom[22796] = 8'he4 ;
            rom[22797] = 8'hff ;
            rom[22798] = 8'hfe ;
            rom[22799] = 8'h1c ;
            rom[22800] = 8'he9 ;
            rom[22801] = 8'hf1 ;
            rom[22802] = 8'h2b ;
            rom[22803] = 8'hfb ;
            rom[22804] = 8'h07 ;
            rom[22805] = 8'hf8 ;
            rom[22806] = 8'hee ;
            rom[22807] = 8'hfa ;
            rom[22808] = 8'hd7 ;
            rom[22809] = 8'h37 ;
            rom[22810] = 8'hf9 ;
            rom[22811] = 8'hef ;
            rom[22812] = 8'h00 ;
            rom[22813] = 8'h13 ;
            rom[22814] = 8'h09 ;
            rom[22815] = 8'hf4 ;
            rom[22816] = 8'heb ;
            rom[22817] = 8'hff ;
            rom[22818] = 8'h1a ;
            rom[22819] = 8'hde ;
            rom[22820] = 8'hfc ;
            rom[22821] = 8'hfb ;
            rom[22822] = 8'hdf ;
            rom[22823] = 8'hfe ;
            rom[22824] = 8'h28 ;
            rom[22825] = 8'h3b ;
            rom[22826] = 8'hff ;
            rom[22827] = 8'h08 ;
            rom[22828] = 8'hfe ;
            rom[22829] = 8'h1c ;
            rom[22830] = 8'h09 ;
            rom[22831] = 8'h1a ;
            rom[22832] = 8'hf9 ;
            rom[22833] = 8'hc0 ;
            rom[22834] = 8'h21 ;
            rom[22835] = 8'h08 ;
            rom[22836] = 8'hfa ;
            rom[22837] = 8'h24 ;
            rom[22838] = 8'he1 ;
            rom[22839] = 8'h0f ;
            rom[22840] = 8'he9 ;
            rom[22841] = 8'hf4 ;
            rom[22842] = 8'hfe ;
            rom[22843] = 8'hfc ;
            rom[22844] = 8'h18 ;
            rom[22845] = 8'hd8 ;
            rom[22846] = 8'h08 ;
            rom[22847] = 8'h1a ;
            rom[22848] = 8'he3 ;
            rom[22849] = 8'h0e ;
            rom[22850] = 8'h13 ;
            rom[22851] = 8'hfe ;
            rom[22852] = 8'hec ;
            rom[22853] = 8'h04 ;
            rom[22854] = 8'hff ;
            rom[22855] = 8'hef ;
            rom[22856] = 8'hd9 ;
            rom[22857] = 8'h03 ;
            rom[22858] = 8'h19 ;
            rom[22859] = 8'h17 ;
            rom[22860] = 8'h0a ;
            rom[22861] = 8'h08 ;
            rom[22862] = 8'he1 ;
            rom[22863] = 8'h0e ;
            rom[22864] = 8'h09 ;
            rom[22865] = 8'h0a ;
            rom[22866] = 8'h03 ;
            rom[22867] = 8'hec ;
            rom[22868] = 8'he8 ;
            rom[22869] = 8'h01 ;
            rom[22870] = 8'hfa ;
            rom[22871] = 8'h36 ;
            rom[22872] = 8'hc9 ;
            rom[22873] = 8'hfd ;
            rom[22874] = 8'h09 ;
            rom[22875] = 8'hfb ;
            rom[22876] = 8'hdd ;
            rom[22877] = 8'hcf ;
            rom[22878] = 8'h20 ;
            rom[22879] = 8'h01 ;
            rom[22880] = 8'h0d ;
            rom[22881] = 8'h2e ;
            rom[22882] = 8'hd2 ;
            rom[22883] = 8'hf9 ;
            rom[22884] = 8'hb1 ;
            rom[22885] = 8'hfb ;
            rom[22886] = 8'hfd ;
            rom[22887] = 8'h04 ;
            rom[22888] = 8'hef ;
            rom[22889] = 8'h0d ;
            rom[22890] = 8'h1f ;
            rom[22891] = 8'hd2 ;
            rom[22892] = 8'h01 ;
            rom[22893] = 8'hd7 ;
            rom[22894] = 8'h05 ;
            rom[22895] = 8'he7 ;
            rom[22896] = 8'hfd ;
            rom[22897] = 8'hfa ;
            rom[22898] = 8'h02 ;
            rom[22899] = 8'h0c ;
            rom[22900] = 8'h1d ;
            rom[22901] = 8'h17 ;
            rom[22902] = 8'h01 ;
            rom[22903] = 8'hee ;
            rom[22904] = 8'h31 ;
            rom[22905] = 8'hc9 ;
            rom[22906] = 8'h11 ;
            rom[22907] = 8'h00 ;
            rom[22908] = 8'h0d ;
            rom[22909] = 8'h07 ;
            rom[22910] = 8'h15 ;
            rom[22911] = 8'he6 ;
            rom[22912] = 8'hf0 ;
            rom[22913] = 8'hf1 ;
            rom[22914] = 8'hf4 ;
            rom[22915] = 8'hed ;
            rom[22916] = 8'h07 ;
            rom[22917] = 8'h28 ;
            rom[22918] = 8'hfb ;
            rom[22919] = 8'h0c ;
            rom[22920] = 8'h49 ;
            rom[22921] = 8'hd8 ;
            rom[22922] = 8'h1c ;
            rom[22923] = 8'hef ;
            rom[22924] = 8'h1e ;
            rom[22925] = 8'h13 ;
            rom[22926] = 8'hf1 ;
            rom[22927] = 8'hce ;
            rom[22928] = 8'hbf ;
            rom[22929] = 8'h1d ;
            rom[22930] = 8'h0c ;
            rom[22931] = 8'h0f ;
            rom[22932] = 8'hed ;
            rom[22933] = 8'hda ;
            rom[22934] = 8'hf2 ;
            rom[22935] = 8'h18 ;
            rom[22936] = 8'hf6 ;
            rom[22937] = 8'hfe ;
            rom[22938] = 8'hd3 ;
            rom[22939] = 8'h10 ;
            rom[22940] = 8'h10 ;
            rom[22941] = 8'h05 ;
            rom[22942] = 8'h0a ;
            rom[22943] = 8'h0c ;
            rom[22944] = 8'hd8 ;
            rom[22945] = 8'hd4 ;
            rom[22946] = 8'hfa ;
            rom[22947] = 8'h1e ;
            rom[22948] = 8'hfc ;
            rom[22949] = 8'hda ;
            rom[22950] = 8'h2d ;
            rom[22951] = 8'hf6 ;
            rom[22952] = 8'hed ;
            rom[22953] = 8'hdf ;
            rom[22954] = 8'h1e ;
            rom[22955] = 8'h1e ;
            rom[22956] = 8'hca ;
            rom[22957] = 8'he5 ;
            rom[22958] = 8'h13 ;
            rom[22959] = 8'hb8 ;
            rom[22960] = 8'h14 ;
            rom[22961] = 8'heb ;
            rom[22962] = 8'hf4 ;
            rom[22963] = 8'hef ;
            rom[22964] = 8'h09 ;
            rom[22965] = 8'hcb ;
            rom[22966] = 8'hf6 ;
            rom[22967] = 8'h26 ;
            rom[22968] = 8'h03 ;
            rom[22969] = 8'hef ;
            rom[22970] = 8'h06 ;
            rom[22971] = 8'hf5 ;
            rom[22972] = 8'hff ;
            rom[22973] = 8'hea ;
            rom[22974] = 8'hfa ;
            rom[22975] = 8'hfc ;
            rom[22976] = 8'hf4 ;
            rom[22977] = 8'hf1 ;
            rom[22978] = 8'h02 ;
            rom[22979] = 8'he9 ;
            rom[22980] = 8'hea ;
            rom[22981] = 8'hf7 ;
            rom[22982] = 8'h1b ;
            rom[22983] = 8'he3 ;
            rom[22984] = 8'h0d ;
            rom[22985] = 8'hfc ;
            rom[22986] = 8'hed ;
            rom[22987] = 8'he4 ;
            rom[22988] = 8'h02 ;
            rom[22989] = 8'h02 ;
            rom[22990] = 8'h02 ;
            rom[22991] = 8'he8 ;
            rom[22992] = 8'h04 ;
            rom[22993] = 8'h0e ;
            rom[22994] = 8'hf3 ;
            rom[22995] = 8'h04 ;
            rom[22996] = 8'hf8 ;
            rom[22997] = 8'h13 ;
            rom[22998] = 8'he3 ;
            rom[22999] = 8'hf2 ;
            rom[23000] = 8'he3 ;
            rom[23001] = 8'hdf ;
            rom[23002] = 8'hbf ;
            rom[23003] = 8'h1e ;
            rom[23004] = 8'h05 ;
            rom[23005] = 8'h0f ;
            rom[23006] = 8'he6 ;
            rom[23007] = 8'hee ;
            rom[23008] = 8'h1d ;
            rom[23009] = 8'he6 ;
            rom[23010] = 8'h05 ;
            rom[23011] = 8'h0a ;
            rom[23012] = 8'h15 ;
            rom[23013] = 8'h16 ;
            rom[23014] = 8'hfd ;
            rom[23015] = 8'h17 ;
            rom[23016] = 8'hf3 ;
            rom[23017] = 8'he7 ;
            rom[23018] = 8'h04 ;
            rom[23019] = 8'h18 ;
            rom[23020] = 8'h1c ;
            rom[23021] = 8'hbd ;
            rom[23022] = 8'h0c ;
            rom[23023] = 8'hed ;
            rom[23024] = 8'hd0 ;
            rom[23025] = 8'h15 ;
            rom[23026] = 8'h1c ;
            rom[23027] = 8'h28 ;
            rom[23028] = 8'h1b ;
            rom[23029] = 8'h09 ;
            rom[23030] = 8'he8 ;
            rom[23031] = 8'hf0 ;
            rom[23032] = 8'he5 ;
            rom[23033] = 8'he6 ;
            rom[23034] = 8'h07 ;
            rom[23035] = 8'h17 ;
            rom[23036] = 8'hfb ;
            rom[23037] = 8'he6 ;
            rom[23038] = 8'h1b ;
            rom[23039] = 8'hf5 ;
            rom[23040] = 8'hf3 ;
            rom[23041] = 8'h23 ;
            rom[23042] = 8'h0d ;
            rom[23043] = 8'h0e ;
            rom[23044] = 8'h03 ;
            rom[23045] = 8'hff ;
            rom[23046] = 8'hf8 ;
            rom[23047] = 8'hd4 ;
            rom[23048] = 8'he6 ;
            rom[23049] = 8'h01 ;
            rom[23050] = 8'h35 ;
            rom[23051] = 8'h0f ;
            rom[23052] = 8'hee ;
            rom[23053] = 8'hfc ;
            rom[23054] = 8'hd7 ;
            rom[23055] = 8'h04 ;
            rom[23056] = 8'h19 ;
            rom[23057] = 8'hf4 ;
            rom[23058] = 8'he3 ;
            rom[23059] = 8'he1 ;
            rom[23060] = 8'h10 ;
            rom[23061] = 8'hf8 ;
            rom[23062] = 8'h15 ;
            rom[23063] = 8'hce ;
            rom[23064] = 8'h01 ;
            rom[23065] = 8'h0d ;
            rom[23066] = 8'he9 ;
            rom[23067] = 8'he7 ;
            rom[23068] = 8'h01 ;
            rom[23069] = 8'hce ;
            rom[23070] = 8'heb ;
            rom[23071] = 8'hf7 ;
            rom[23072] = 8'hfc ;
            rom[23073] = 8'h27 ;
            rom[23074] = 8'hef ;
            rom[23075] = 8'he6 ;
            rom[23076] = 8'hf2 ;
            rom[23077] = 8'hf6 ;
            rom[23078] = 8'he8 ;
            rom[23079] = 8'h0d ;
            rom[23080] = 8'hf1 ;
            rom[23081] = 8'hf0 ;
            rom[23082] = 8'h24 ;
            rom[23083] = 8'h06 ;
            rom[23084] = 8'hf0 ;
            rom[23085] = 8'hea ;
            rom[23086] = 8'hf7 ;
            rom[23087] = 8'hf8 ;
            rom[23088] = 8'hef ;
            rom[23089] = 8'hf6 ;
            rom[23090] = 8'he9 ;
            rom[23091] = 8'hf1 ;
            rom[23092] = 8'hd8 ;
            rom[23093] = 8'h06 ;
            rom[23094] = 8'heb ;
            rom[23095] = 8'h12 ;
            rom[23096] = 8'hf5 ;
            rom[23097] = 8'hfd ;
            rom[23098] = 8'heb ;
            rom[23099] = 8'h0b ;
            rom[23100] = 8'h13 ;
            rom[23101] = 8'h0b ;
            rom[23102] = 8'h14 ;
            rom[23103] = 8'h03 ;
            rom[23104] = 8'hed ;
            rom[23105] = 8'h06 ;
            rom[23106] = 8'h07 ;
            rom[23107] = 8'hf2 ;
            rom[23108] = 8'hd1 ;
            rom[23109] = 8'h08 ;
            rom[23110] = 8'hec ;
            rom[23111] = 8'hfd ;
            rom[23112] = 8'hf0 ;
            rom[23113] = 8'hd6 ;
            rom[23114] = 8'h11 ;
            rom[23115] = 8'he9 ;
            rom[23116] = 8'hb6 ;
            rom[23117] = 8'hc4 ;
            rom[23118] = 8'he9 ;
            rom[23119] = 8'hd7 ;
            rom[23120] = 8'hf5 ;
            rom[23121] = 8'hea ;
            rom[23122] = 8'he8 ;
            rom[23123] = 8'hd5 ;
            rom[23124] = 8'he9 ;
            rom[23125] = 8'hdb ;
            rom[23126] = 8'h08 ;
            rom[23127] = 8'hfd ;
            rom[23128] = 8'he6 ;
            rom[23129] = 8'hfe ;
            rom[23130] = 8'hf3 ;
            rom[23131] = 8'hf5 ;
            rom[23132] = 8'hed ;
            rom[23133] = 8'hfa ;
            rom[23134] = 8'hee ;
            rom[23135] = 8'he5 ;
            rom[23136] = 8'hd4 ;
            rom[23137] = 8'h1d ;
            rom[23138] = 8'hee ;
            rom[23139] = 8'hf4 ;
            rom[23140] = 8'hef ;
            rom[23141] = 8'h0c ;
            rom[23142] = 8'h11 ;
            rom[23143] = 8'h09 ;
            rom[23144] = 8'hed ;
            rom[23145] = 8'h0e ;
            rom[23146] = 8'hed ;
            rom[23147] = 8'hfc ;
            rom[23148] = 8'h10 ;
            rom[23149] = 8'hef ;
            rom[23150] = 8'hfc ;
            rom[23151] = 8'h09 ;
            rom[23152] = 8'h04 ;
            rom[23153] = 8'h05 ;
            rom[23154] = 8'h1b ;
            rom[23155] = 8'h04 ;
            rom[23156] = 8'hf3 ;
            rom[23157] = 8'h1a ;
            rom[23158] = 8'h1c ;
            rom[23159] = 8'h07 ;
            rom[23160] = 8'hfd ;
            rom[23161] = 8'hf1 ;
            rom[23162] = 8'h0c ;
            rom[23163] = 8'hf0 ;
            rom[23164] = 8'hc7 ;
            rom[23165] = 8'h2b ;
            rom[23166] = 8'h06 ;
            rom[23167] = 8'h02 ;
            rom[23168] = 8'hde ;
            rom[23169] = 8'h17 ;
            rom[23170] = 8'h15 ;
            rom[23171] = 8'h14 ;
            rom[23172] = 8'h31 ;
            rom[23173] = 8'h0e ;
            rom[23174] = 8'hfd ;
            rom[23175] = 8'h1f ;
            rom[23176] = 8'h03 ;
            rom[23177] = 8'h15 ;
            rom[23178] = 8'hf1 ;
            rom[23179] = 8'hf1 ;
            rom[23180] = 8'hf2 ;
            rom[23181] = 8'h32 ;
            rom[23182] = 8'h13 ;
            rom[23183] = 8'h10 ;
            rom[23184] = 8'h12 ;
            rom[23185] = 8'h1a ;
            rom[23186] = 8'hf8 ;
            rom[23187] = 8'hce ;
            rom[23188] = 8'h07 ;
            rom[23189] = 8'hf0 ;
            rom[23190] = 8'h1d ;
            rom[23191] = 8'h02 ;
            rom[23192] = 8'he3 ;
            rom[23193] = 8'hf8 ;
            rom[23194] = 8'h03 ;
            rom[23195] = 8'h0a ;
            rom[23196] = 8'h04 ;
            rom[23197] = 8'hf8 ;
            rom[23198] = 8'hf4 ;
            rom[23199] = 8'h1f ;
            rom[23200] = 8'h32 ;
            rom[23201] = 8'hf2 ;
            rom[23202] = 8'h14 ;
            rom[23203] = 8'hc8 ;
            rom[23204] = 8'hc2 ;
            rom[23205] = 8'hf9 ;
            rom[23206] = 8'h2f ;
            rom[23207] = 8'hf5 ;
            rom[23208] = 8'h0d ;
            rom[23209] = 8'h0a ;
            rom[23210] = 8'hd4 ;
            rom[23211] = 8'h13 ;
            rom[23212] = 8'hff ;
            rom[23213] = 8'h05 ;
            rom[23214] = 8'hf2 ;
            rom[23215] = 8'h21 ;
            rom[23216] = 8'he4 ;
            rom[23217] = 8'hf2 ;
            rom[23218] = 8'he2 ;
            rom[23219] = 8'hf3 ;
            rom[23220] = 8'hf4 ;
            rom[23221] = 8'hdf ;
            rom[23222] = 8'hf1 ;
            rom[23223] = 8'hf0 ;
            rom[23224] = 8'heb ;
            rom[23225] = 8'hd3 ;
            rom[23226] = 8'hc5 ;
            rom[23227] = 8'h00 ;
            rom[23228] = 8'hf1 ;
            rom[23229] = 8'h01 ;
            rom[23230] = 8'hf9 ;
            rom[23231] = 8'h18 ;
            rom[23232] = 8'h3c ;
            rom[23233] = 8'hfc ;
            rom[23234] = 8'h06 ;
            rom[23235] = 8'h1f ;
            rom[23236] = 8'h08 ;
            rom[23237] = 8'h13 ;
            rom[23238] = 8'h0c ;
            rom[23239] = 8'hff ;
            rom[23240] = 8'he5 ;
            rom[23241] = 8'hf2 ;
            rom[23242] = 8'hdb ;
            rom[23243] = 8'hea ;
            rom[23244] = 8'h1d ;
            rom[23245] = 8'hd8 ;
            rom[23246] = 8'hc6 ;
            rom[23247] = 8'h1a ;
            rom[23248] = 8'hf5 ;
            rom[23249] = 8'he8 ;
            rom[23250] = 8'h1a ;
            rom[23251] = 8'h1b ;
            rom[23252] = 8'hf6 ;
            rom[23253] = 8'h00 ;
            rom[23254] = 8'hef ;
            rom[23255] = 8'h09 ;
            rom[23256] = 8'he2 ;
            rom[23257] = 8'hce ;
            rom[23258] = 8'hf8 ;
            rom[23259] = 8'h1e ;
            rom[23260] = 8'h1b ;
            rom[23261] = 8'h1f ;
            rom[23262] = 8'h0d ;
            rom[23263] = 8'h0e ;
            rom[23264] = 8'h07 ;
            rom[23265] = 8'h2c ;
            rom[23266] = 8'hd4 ;
            rom[23267] = 8'h05 ;
            rom[23268] = 8'he4 ;
            rom[23269] = 8'h1f ;
            rom[23270] = 8'h1d ;
            rom[23271] = 8'hec ;
            rom[23272] = 8'hfc ;
            rom[23273] = 8'h0d ;
            rom[23274] = 8'h2a ;
            rom[23275] = 8'hef ;
            rom[23276] = 8'hdf ;
            rom[23277] = 8'h01 ;
            rom[23278] = 8'hcc ;
            rom[23279] = 8'hfa ;
            rom[23280] = 8'h30 ;
            rom[23281] = 8'h08 ;
            rom[23282] = 8'h11 ;
            rom[23283] = 8'h23 ;
            rom[23284] = 8'he3 ;
            rom[23285] = 8'he8 ;
            rom[23286] = 8'hdf ;
            rom[23287] = 8'h09 ;
            rom[23288] = 8'hc1 ;
            rom[23289] = 8'h13 ;
            rom[23290] = 8'hee ;
            rom[23291] = 8'hf9 ;
            rom[23292] = 8'h03 ;
            rom[23293] = 8'h20 ;
            rom[23294] = 8'h20 ;
            rom[23295] = 8'hff ;
            rom[23296] = 8'h0a ;
            rom[23297] = 8'hbd ;
            rom[23298] = 8'hcd ;
            rom[23299] = 8'h0b ;
            rom[23300] = 8'hf4 ;
            rom[23301] = 8'h24 ;
            rom[23302] = 8'hea ;
            rom[23303] = 8'hec ;
            rom[23304] = 8'hfc ;
            rom[23305] = 8'he4 ;
            rom[23306] = 8'hdf ;
            rom[23307] = 8'hf8 ;
            rom[23308] = 8'he1 ;
            rom[23309] = 8'h0c ;
            rom[23310] = 8'h10 ;
            rom[23311] = 8'hf3 ;
            rom[23312] = 8'h03 ;
            rom[23313] = 8'hff ;
            rom[23314] = 8'h07 ;
            rom[23315] = 8'hfa ;
            rom[23316] = 8'h0b ;
            rom[23317] = 8'h07 ;
            rom[23318] = 8'hee ;
            rom[23319] = 8'h08 ;
            rom[23320] = 8'hd6 ;
            rom[23321] = 8'h18 ;
            rom[23322] = 8'he8 ;
            rom[23323] = 8'hf0 ;
            rom[23324] = 8'he4 ;
            rom[23325] = 8'h0a ;
            rom[23326] = 8'h01 ;
            rom[23327] = 8'h0d ;
            rom[23328] = 8'hc5 ;
            rom[23329] = 8'hcf ;
            rom[23330] = 8'hf3 ;
            rom[23331] = 8'h0b ;
            rom[23332] = 8'hd1 ;
            rom[23333] = 8'hb9 ;
            rom[23334] = 8'h02 ;
            rom[23335] = 8'hf5 ;
            rom[23336] = 8'hea ;
            rom[23337] = 8'hf8 ;
            rom[23338] = 8'h11 ;
            rom[23339] = 8'h0e ;
            rom[23340] = 8'he3 ;
            rom[23341] = 8'hf1 ;
            rom[23342] = 8'he2 ;
            rom[23343] = 8'h1a ;
            rom[23344] = 8'hfc ;
            rom[23345] = 8'hcf ;
            rom[23346] = 8'hff ;
            rom[23347] = 8'h03 ;
            rom[23348] = 8'h12 ;
            rom[23349] = 8'he5 ;
            rom[23350] = 8'h1b ;
            rom[23351] = 8'h26 ;
            rom[23352] = 8'he8 ;
            rom[23353] = 8'hfd ;
            rom[23354] = 8'hfb ;
            rom[23355] = 8'hf3 ;
            rom[23356] = 8'hd4 ;
            rom[23357] = 8'hea ;
            rom[23358] = 8'h0c ;
            rom[23359] = 8'h0c ;
            rom[23360] = 8'hf0 ;
            rom[23361] = 8'h14 ;
            rom[23362] = 8'hef ;
            rom[23363] = 8'h02 ;
            rom[23364] = 8'h17 ;
            rom[23365] = 8'hf0 ;
            rom[23366] = 8'hfe ;
            rom[23367] = 8'hf7 ;
            rom[23368] = 8'h1c ;
            rom[23369] = 8'hff ;
            rom[23370] = 8'h07 ;
            rom[23371] = 8'hf5 ;
            rom[23372] = 8'h30 ;
            rom[23373] = 8'hdb ;
            rom[23374] = 8'hf8 ;
            rom[23375] = 8'h1f ;
            rom[23376] = 8'h17 ;
            rom[23377] = 8'h29 ;
            rom[23378] = 8'h0f ;
            rom[23379] = 8'hfd ;
            rom[23380] = 8'hf6 ;
            rom[23381] = 8'h12 ;
            rom[23382] = 8'hfa ;
            rom[23383] = 8'he3 ;
            rom[23384] = 8'h1c ;
            rom[23385] = 8'hd5 ;
            rom[23386] = 8'h0b ;
            rom[23387] = 8'hfe ;
            rom[23388] = 8'h03 ;
            rom[23389] = 8'hec ;
            rom[23390] = 8'hfa ;
            rom[23391] = 8'h11 ;
            rom[23392] = 8'h14 ;
            rom[23393] = 8'hfa ;
            rom[23394] = 8'h07 ;
            rom[23395] = 8'he9 ;
            rom[23396] = 8'hf7 ;
            rom[23397] = 8'hda ;
            rom[23398] = 8'h01 ;
            rom[23399] = 8'h0d ;
            rom[23400] = 8'hee ;
            rom[23401] = 8'hed ;
            rom[23402] = 8'h0a ;
            rom[23403] = 8'h13 ;
            rom[23404] = 8'h01 ;
            rom[23405] = 8'hf7 ;
            rom[23406] = 8'h18 ;
            rom[23407] = 8'hed ;
            rom[23408] = 8'hca ;
            rom[23409] = 8'h0c ;
            rom[23410] = 8'h02 ;
            rom[23411] = 8'hed ;
            rom[23412] = 8'h00 ;
            rom[23413] = 8'hea ;
            rom[23414] = 8'he0 ;
            rom[23415] = 8'h15 ;
            rom[23416] = 8'h11 ;
            rom[23417] = 8'he6 ;
            rom[23418] = 8'hf2 ;
            rom[23419] = 8'hf0 ;
            rom[23420] = 8'hff ;
            rom[23421] = 8'h06 ;
            rom[23422] = 8'h23 ;
            rom[23423] = 8'he8 ;
            rom[23424] = 8'hfe ;
            rom[23425] = 8'hc8 ;
            rom[23426] = 8'hdd ;
            rom[23427] = 8'h0f ;
            rom[23428] = 8'h0c ;
            rom[23429] = 8'hbe ;
            rom[23430] = 8'he5 ;
            rom[23431] = 8'he5 ;
            rom[23432] = 8'heb ;
            rom[23433] = 8'h13 ;
            rom[23434] = 8'h0d ;
            rom[23435] = 8'h00 ;
            rom[23436] = 8'he0 ;
            rom[23437] = 8'hff ;
            rom[23438] = 8'hf9 ;
            rom[23439] = 8'hf4 ;
            rom[23440] = 8'hf7 ;
            rom[23441] = 8'hdd ;
            rom[23442] = 8'hed ;
            rom[23443] = 8'hef ;
            rom[23444] = 8'h22 ;
            rom[23445] = 8'h18 ;
            rom[23446] = 8'he0 ;
            rom[23447] = 8'h05 ;
            rom[23448] = 8'hc0 ;
            rom[23449] = 8'h17 ;
            rom[23450] = 8'hea ;
            rom[23451] = 8'hc5 ;
            rom[23452] = 8'h16 ;
            rom[23453] = 8'hf8 ;
            rom[23454] = 8'hf4 ;
            rom[23455] = 8'h0e ;
            rom[23456] = 8'hfb ;
            rom[23457] = 8'hf5 ;
            rom[23458] = 8'h12 ;
            rom[23459] = 8'hd2 ;
            rom[23460] = 8'hf8 ;
            rom[23461] = 8'hd9 ;
            rom[23462] = 8'h05 ;
            rom[23463] = 8'h08 ;
            rom[23464] = 8'h2c ;
            rom[23465] = 8'he7 ;
            rom[23466] = 8'hc4 ;
            rom[23467] = 8'hd2 ;
            rom[23468] = 8'h05 ;
            rom[23469] = 8'hf3 ;
            rom[23470] = 8'hf4 ;
            rom[23471] = 8'hf7 ;
            rom[23472] = 8'hcd ;
            rom[23473] = 8'hf9 ;
            rom[23474] = 8'hf8 ;
            rom[23475] = 8'h00 ;
            rom[23476] = 8'he8 ;
            rom[23477] = 8'hf7 ;
            rom[23478] = 8'hd6 ;
            rom[23479] = 8'hc5 ;
            rom[23480] = 8'hfe ;
            rom[23481] = 8'h08 ;
            rom[23482] = 8'he7 ;
            rom[23483] = 8'hf7 ;
            rom[23484] = 8'h12 ;
            rom[23485] = 8'h11 ;
            rom[23486] = 8'h05 ;
            rom[23487] = 8'he6 ;
            rom[23488] = 8'hda ;
            rom[23489] = 8'hf6 ;
            rom[23490] = 8'h11 ;
            rom[23491] = 8'he8 ;
            rom[23492] = 8'h1e ;
            rom[23493] = 8'hf3 ;
            rom[23494] = 8'hcd ;
            rom[23495] = 8'hf4 ;
            rom[23496] = 8'hdf ;
            rom[23497] = 8'h0f ;
            rom[23498] = 8'h22 ;
            rom[23499] = 8'h1f ;
            rom[23500] = 8'h00 ;
            rom[23501] = 8'hf4 ;
            rom[23502] = 8'hf0 ;
            rom[23503] = 8'h0c ;
            rom[23504] = 8'hd4 ;
            rom[23505] = 8'hee ;
            rom[23506] = 8'hd9 ;
            rom[23507] = 8'hc9 ;
            rom[23508] = 8'hde ;
            rom[23509] = 8'h1d ;
            rom[23510] = 8'h05 ;
            rom[23511] = 8'hf6 ;
            rom[23512] = 8'hf5 ;
            rom[23513] = 8'hf7 ;
            rom[23514] = 8'h31 ;
            rom[23515] = 8'h16 ;
            rom[23516] = 8'he4 ;
            rom[23517] = 8'hfa ;
            rom[23518] = 8'h00 ;
            rom[23519] = 8'h01 ;
            rom[23520] = 8'h12 ;
            rom[23521] = 8'h10 ;
            rom[23522] = 8'h25 ;
            rom[23523] = 8'he6 ;
            rom[23524] = 8'hd7 ;
            rom[23525] = 8'hf2 ;
            rom[23526] = 8'heb ;
            rom[23527] = 8'hda ;
            rom[23528] = 8'he5 ;
            rom[23529] = 8'h05 ;
            rom[23530] = 8'h2b ;
            rom[23531] = 8'h05 ;
            rom[23532] = 8'hff ;
            rom[23533] = 8'hfb ;
            rom[23534] = 8'hec ;
            rom[23535] = 8'he7 ;
            rom[23536] = 8'he1 ;
            rom[23537] = 8'hfb ;
            rom[23538] = 8'h16 ;
            rom[23539] = 8'h0a ;
            rom[23540] = 8'hef ;
            rom[23541] = 8'h06 ;
            rom[23542] = 8'hfc ;
            rom[23543] = 8'hf3 ;
            rom[23544] = 8'hf2 ;
            rom[23545] = 8'hfd ;
            rom[23546] = 8'hc0 ;
            rom[23547] = 8'hed ;
            rom[23548] = 8'h09 ;
            rom[23549] = 8'h06 ;
            rom[23550] = 8'hf4 ;
            rom[23551] = 8'hd4 ;
            rom[23552] = 8'h01 ;
            rom[23553] = 8'h0e ;
            rom[23554] = 8'he8 ;
            rom[23555] = 8'hfc ;
            rom[23556] = 8'h1d ;
            rom[23557] = 8'he4 ;
            rom[23558] = 8'hf2 ;
            rom[23559] = 8'he7 ;
            rom[23560] = 8'hdd ;
            rom[23561] = 8'hf5 ;
            rom[23562] = 8'hed ;
            rom[23563] = 8'h0e ;
            rom[23564] = 8'h11 ;
            rom[23565] = 8'hf9 ;
            rom[23566] = 8'h0b ;
            rom[23567] = 8'hfd ;
            rom[23568] = 8'hb3 ;
            rom[23569] = 8'hdb ;
            rom[23570] = 8'h09 ;
            rom[23571] = 8'hd3 ;
            rom[23572] = 8'h02 ;
            rom[23573] = 8'hf6 ;
            rom[23574] = 8'he9 ;
            rom[23575] = 8'hdd ;
            rom[23576] = 8'hc7 ;
            rom[23577] = 8'h03 ;
            rom[23578] = 8'hef ;
            rom[23579] = 8'h08 ;
            rom[23580] = 8'he4 ;
            rom[23581] = 8'hcb ;
            rom[23582] = 8'hf3 ;
            rom[23583] = 8'h0b ;
            rom[23584] = 8'hf8 ;
            rom[23585] = 8'hf3 ;
            rom[23586] = 8'hc7 ;
            rom[23587] = 8'hbb ;
            rom[23588] = 8'h0d ;
            rom[23589] = 8'hee ;
            rom[23590] = 8'h19 ;
            rom[23591] = 8'h01 ;
            rom[23592] = 8'h2a ;
            rom[23593] = 8'h08 ;
            rom[23594] = 8'h10 ;
            rom[23595] = 8'he6 ;
            rom[23596] = 8'hfb ;
            rom[23597] = 8'h05 ;
            rom[23598] = 8'h02 ;
            rom[23599] = 8'he6 ;
            rom[23600] = 8'h00 ;
            rom[23601] = 8'he0 ;
            rom[23602] = 8'hea ;
            rom[23603] = 8'h0d ;
            rom[23604] = 8'h16 ;
            rom[23605] = 8'hf6 ;
            rom[23606] = 8'h1c ;
            rom[23607] = 8'hc8 ;
            rom[23608] = 8'hec ;
            rom[23609] = 8'he6 ;
            rom[23610] = 8'hff ;
            rom[23611] = 8'hfc ;
            rom[23612] = 8'h04 ;
            rom[23613] = 8'h18 ;
            rom[23614] = 8'he8 ;
            rom[23615] = 8'h03 ;
            rom[23616] = 8'h06 ;
            rom[23617] = 8'hce ;
            rom[23618] = 8'h0c ;
            rom[23619] = 8'h00 ;
            rom[23620] = 8'hfc ;
            rom[23621] = 8'hf9 ;
            rom[23622] = 8'hfc ;
            rom[23623] = 8'h0f ;
            rom[23624] = 8'hfb ;
            rom[23625] = 8'hd9 ;
            rom[23626] = 8'hea ;
            rom[23627] = 8'h1f ;
            rom[23628] = 8'hd4 ;
            rom[23629] = 8'he6 ;
            rom[23630] = 8'he9 ;
            rom[23631] = 8'hf0 ;
            rom[23632] = 8'hd2 ;
            rom[23633] = 8'hd2 ;
            rom[23634] = 8'hde ;
            rom[23635] = 8'he9 ;
            rom[23636] = 8'hed ;
            rom[23637] = 8'hf1 ;
            rom[23638] = 8'hf5 ;
            rom[23639] = 8'h0d ;
            rom[23640] = 8'h08 ;
            rom[23641] = 8'hf9 ;
            rom[23642] = 8'hfc ;
            rom[23643] = 8'h10 ;
            rom[23644] = 8'hd0 ;
            rom[23645] = 8'he5 ;
            rom[23646] = 8'hf8 ;
            rom[23647] = 8'hd6 ;
            rom[23648] = 8'he7 ;
            rom[23649] = 8'h06 ;
            rom[23650] = 8'hee ;
            rom[23651] = 8'hdd ;
            rom[23652] = 8'hf6 ;
            rom[23653] = 8'h0d ;
            rom[23654] = 8'h31 ;
            rom[23655] = 8'hf7 ;
            rom[23656] = 8'hf2 ;
            rom[23657] = 8'hf7 ;
            rom[23658] = 8'he5 ;
            rom[23659] = 8'hef ;
            rom[23660] = 8'hf6 ;
            rom[23661] = 8'h0b ;
            rom[23662] = 8'hd8 ;
            rom[23663] = 8'h33 ;
            rom[23664] = 8'h19 ;
            rom[23665] = 8'h1b ;
            rom[23666] = 8'h25 ;
            rom[23667] = 8'hf7 ;
            rom[23668] = 8'hea ;
            rom[23669] = 8'h08 ;
            rom[23670] = 8'hfd ;
            rom[23671] = 8'hf7 ;
            rom[23672] = 8'h11 ;
            rom[23673] = 8'h08 ;
            rom[23674] = 8'hff ;
            rom[23675] = 8'h17 ;
            rom[23676] = 8'h26 ;
            rom[23677] = 8'hf9 ;
            rom[23678] = 8'h01 ;
            rom[23679] = 8'he4 ;
            rom[23680] = 8'h1d ;
            rom[23681] = 8'hd5 ;
            rom[23682] = 8'h01 ;
            rom[23683] = 8'h03 ;
            rom[23684] = 8'hfc ;
            rom[23685] = 8'h0b ;
            rom[23686] = 8'h09 ;
            rom[23687] = 8'h05 ;
            rom[23688] = 8'h26 ;
            rom[23689] = 8'hda ;
            rom[23690] = 8'hfe ;
            rom[23691] = 8'hd3 ;
            rom[23692] = 8'hef ;
            rom[23693] = 8'he1 ;
            rom[23694] = 8'hf1 ;
            rom[23695] = 8'hf0 ;
            rom[23696] = 8'hdb ;
            rom[23697] = 8'he8 ;
            rom[23698] = 8'h03 ;
            rom[23699] = 8'h01 ;
            rom[23700] = 8'h0e ;
            rom[23701] = 8'hcd ;
            rom[23702] = 8'hbf ;
            rom[23703] = 8'h2c ;
            rom[23704] = 8'h0a ;
            rom[23705] = 8'hfe ;
            rom[23706] = 8'h05 ;
            rom[23707] = 8'h07 ;
            rom[23708] = 8'hf4 ;
            rom[23709] = 8'h04 ;
            rom[23710] = 8'hf7 ;
            rom[23711] = 8'h05 ;
            rom[23712] = 8'hf5 ;
            rom[23713] = 8'hec ;
            rom[23714] = 8'h17 ;
            rom[23715] = 8'h36 ;
            rom[23716] = 8'h1a ;
            rom[23717] = 8'hfa ;
            rom[23718] = 8'h17 ;
            rom[23719] = 8'hf4 ;
            rom[23720] = 8'hc9 ;
            rom[23721] = 8'hea ;
            rom[23722] = 8'hfb ;
            rom[23723] = 8'h0c ;
            rom[23724] = 8'hf6 ;
            rom[23725] = 8'h1f ;
            rom[23726] = 8'h0b ;
            rom[23727] = 8'hd9 ;
            rom[23728] = 8'hdf ;
            rom[23729] = 8'hec ;
            rom[23730] = 8'hfc ;
            rom[23731] = 8'h02 ;
            rom[23732] = 8'h11 ;
            rom[23733] = 8'hf2 ;
            rom[23734] = 8'hde ;
            rom[23735] = 8'hff ;
            rom[23736] = 8'h0e ;
            rom[23737] = 8'h0c ;
            rom[23738] = 8'h01 ;
            rom[23739] = 8'hdc ;
            rom[23740] = 8'h2d ;
            rom[23741] = 8'hd6 ;
            rom[23742] = 8'hf4 ;
            rom[23743] = 8'hfb ;
            rom[23744] = 8'hc7 ;
            rom[23745] = 8'h2c ;
            rom[23746] = 8'h21 ;
            rom[23747] = 8'h36 ;
            rom[23748] = 8'hfe ;
            rom[23749] = 8'h14 ;
            rom[23750] = 8'h08 ;
            rom[23751] = 8'he6 ;
            rom[23752] = 8'h09 ;
            rom[23753] = 8'h00 ;
            rom[23754] = 8'hdd ;
            rom[23755] = 8'hfe ;
            rom[23756] = 8'h23 ;
            rom[23757] = 8'he8 ;
            rom[23758] = 8'h30 ;
            rom[23759] = 8'h04 ;
            rom[23760] = 8'h1a ;
            rom[23761] = 8'he7 ;
            rom[23762] = 8'h0d ;
            rom[23763] = 8'h01 ;
            rom[23764] = 8'he8 ;
            rom[23765] = 8'hff ;
            rom[23766] = 8'hcc ;
            rom[23767] = 8'hfa ;
            rom[23768] = 8'h43 ;
            rom[23769] = 8'hf9 ;
            rom[23770] = 8'hf9 ;
            rom[23771] = 8'h12 ;
            rom[23772] = 8'h10 ;
            rom[23773] = 8'hfe ;
            rom[23774] = 8'h07 ;
            rom[23775] = 8'h15 ;
            rom[23776] = 8'h06 ;
            rom[23777] = 8'he1 ;
            rom[23778] = 8'he9 ;
            rom[23779] = 8'hfc ;
            rom[23780] = 8'he9 ;
            rom[23781] = 8'h20 ;
            rom[23782] = 8'h13 ;
            rom[23783] = 8'h01 ;
            rom[23784] = 8'hef ;
            rom[23785] = 8'hb0 ;
            rom[23786] = 8'h15 ;
            rom[23787] = 8'h09 ;
            rom[23788] = 8'hf5 ;
            rom[23789] = 8'heb ;
            rom[23790] = 8'h1d ;
            rom[23791] = 8'hda ;
            rom[23792] = 8'hd1 ;
            rom[23793] = 8'hd6 ;
            rom[23794] = 8'h1d ;
            rom[23795] = 8'h0e ;
            rom[23796] = 8'h17 ;
            rom[23797] = 8'h09 ;
            rom[23798] = 8'hf6 ;
            rom[23799] = 8'hd7 ;
            rom[23800] = 8'hdc ;
            rom[23801] = 8'hed ;
            rom[23802] = 8'h0e ;
            rom[23803] = 8'h0a ;
            rom[23804] = 8'hf3 ;
            rom[23805] = 8'hf2 ;
            rom[23806] = 8'h0c ;
            rom[23807] = 8'hef ;
            rom[23808] = 8'hff ;
            rom[23809] = 8'h19 ;
            rom[23810] = 8'h05 ;
            rom[23811] = 8'h08 ;
            rom[23812] = 8'h21 ;
            rom[23813] = 8'h04 ;
            rom[23814] = 8'h05 ;
            rom[23815] = 8'hd3 ;
            rom[23816] = 8'hf0 ;
            rom[23817] = 8'hfa ;
            rom[23818] = 8'he7 ;
            rom[23819] = 8'hbf ;
            rom[23820] = 8'h00 ;
            rom[23821] = 8'h06 ;
            rom[23822] = 8'hfc ;
            rom[23823] = 8'h18 ;
            rom[23824] = 8'hd5 ;
            rom[23825] = 8'h04 ;
            rom[23826] = 8'h07 ;
            rom[23827] = 8'hc8 ;
            rom[23828] = 8'hec ;
            rom[23829] = 8'hf5 ;
            rom[23830] = 8'h0b ;
            rom[23831] = 8'h2a ;
            rom[23832] = 8'h08 ;
            rom[23833] = 8'h24 ;
            rom[23834] = 8'hee ;
            rom[23835] = 8'hf3 ;
            rom[23836] = 8'hfb ;
            rom[23837] = 8'h07 ;
            rom[23838] = 8'h11 ;
            rom[23839] = 8'h0c ;
            rom[23840] = 8'hf0 ;
            rom[23841] = 8'hc4 ;
            rom[23842] = 8'hf4 ;
            rom[23843] = 8'he6 ;
            rom[23844] = 8'h18 ;
            rom[23845] = 8'hd0 ;
            rom[23846] = 8'h23 ;
            rom[23847] = 8'h03 ;
            rom[23848] = 8'he2 ;
            rom[23849] = 8'hb4 ;
            rom[23850] = 8'hf8 ;
            rom[23851] = 8'h1f ;
            rom[23852] = 8'hfa ;
            rom[23853] = 8'hd2 ;
            rom[23854] = 8'h1f ;
            rom[23855] = 8'h09 ;
            rom[23856] = 8'h26 ;
            rom[23857] = 8'he3 ;
            rom[23858] = 8'hf7 ;
            rom[23859] = 8'h11 ;
            rom[23860] = 8'hed ;
            rom[23861] = 8'hf7 ;
            rom[23862] = 8'h08 ;
            rom[23863] = 8'h14 ;
            rom[23864] = 8'h13 ;
            rom[23865] = 8'he8 ;
            rom[23866] = 8'h01 ;
            rom[23867] = 8'h15 ;
            rom[23868] = 8'hf8 ;
            rom[23869] = 8'hfc ;
            rom[23870] = 8'h03 ;
            rom[23871] = 8'h10 ;
            rom[23872] = 8'hfe ;
            rom[23873] = 8'h10 ;
            rom[23874] = 8'hf8 ;
            rom[23875] = 8'he2 ;
            rom[23876] = 8'h18 ;
            rom[23877] = 8'he7 ;
            rom[23878] = 8'he2 ;
            rom[23879] = 8'hec ;
            rom[23880] = 8'h0d ;
            rom[23881] = 8'hec ;
            rom[23882] = 8'hcb ;
            rom[23883] = 8'hf1 ;
            rom[23884] = 8'hfc ;
            rom[23885] = 8'hff ;
            rom[23886] = 8'hf5 ;
            rom[23887] = 8'hf9 ;
            rom[23888] = 8'h21 ;
            rom[23889] = 8'h26 ;
            rom[23890] = 8'h02 ;
            rom[23891] = 8'hff ;
            rom[23892] = 8'h05 ;
            rom[23893] = 8'h0d ;
            rom[23894] = 8'hfa ;
            rom[23895] = 8'h03 ;
            rom[23896] = 8'h0b ;
            rom[23897] = 8'hdb ;
            rom[23898] = 8'hec ;
            rom[23899] = 8'hfa ;
            rom[23900] = 8'h27 ;
            rom[23901] = 8'h14 ;
            rom[23902] = 8'hc9 ;
            rom[23903] = 8'hff ;
            rom[23904] = 8'hf6 ;
            rom[23905] = 8'h02 ;
            rom[23906] = 8'he7 ;
            rom[23907] = 8'h0e ;
            rom[23908] = 8'h24 ;
            rom[23909] = 8'h02 ;
            rom[23910] = 8'h08 ;
            rom[23911] = 8'hf1 ;
            rom[23912] = 8'hc0 ;
            rom[23913] = 8'hcf ;
            rom[23914] = 8'h04 ;
            rom[23915] = 8'h2e ;
            rom[23916] = 8'hf1 ;
            rom[23917] = 8'he5 ;
            rom[23918] = 8'h1b ;
            rom[23919] = 8'h05 ;
            rom[23920] = 8'hdb ;
            rom[23921] = 8'h1a ;
            rom[23922] = 8'h07 ;
            rom[23923] = 8'h1d ;
            rom[23924] = 8'h08 ;
            rom[23925] = 8'h0b ;
            rom[23926] = 8'hcb ;
            rom[23927] = 8'hd0 ;
            rom[23928] = 8'hf9 ;
            rom[23929] = 8'h03 ;
            rom[23930] = 8'h07 ;
            rom[23931] = 8'h3f ;
            rom[23932] = 8'h11 ;
            rom[23933] = 8'hed ;
            rom[23934] = 8'h07 ;
            rom[23935] = 8'h02 ;
            rom[23936] = 8'h29 ;
            rom[23937] = 8'h05 ;
            rom[23938] = 8'hff ;
            rom[23939] = 8'hf5 ;
            rom[23940] = 8'h0f ;
            rom[23941] = 8'hbf ;
            rom[23942] = 8'he6 ;
            rom[23943] = 8'h01 ;
            rom[23944] = 8'hf2 ;
            rom[23945] = 8'he6 ;
            rom[23946] = 8'hd5 ;
            rom[23947] = 8'hef ;
            rom[23948] = 8'hd2 ;
            rom[23949] = 8'he5 ;
            rom[23950] = 8'hcf ;
            rom[23951] = 8'h10 ;
            rom[23952] = 8'he2 ;
            rom[23953] = 8'hfd ;
            rom[23954] = 8'hef ;
            rom[23955] = 8'hf7 ;
            rom[23956] = 8'hfc ;
            rom[23957] = 8'hff ;
            rom[23958] = 8'h04 ;
            rom[23959] = 8'hfb ;
            rom[23960] = 8'h0a ;
            rom[23961] = 8'h00 ;
            rom[23962] = 8'hfc ;
            rom[23963] = 8'hfb ;
            rom[23964] = 8'h10 ;
            rom[23965] = 8'h01 ;
            rom[23966] = 8'hea ;
            rom[23967] = 8'h10 ;
            rom[23968] = 8'h11 ;
            rom[23969] = 8'hef ;
            rom[23970] = 8'h25 ;
            rom[23971] = 8'hd1 ;
            rom[23972] = 8'hca ;
            rom[23973] = 8'hd5 ;
            rom[23974] = 8'hff ;
            rom[23975] = 8'he5 ;
            rom[23976] = 8'hf2 ;
            rom[23977] = 8'hf0 ;
            rom[23978] = 8'he6 ;
            rom[23979] = 8'he4 ;
            rom[23980] = 8'hed ;
            rom[23981] = 8'hee ;
            rom[23982] = 8'hf9 ;
            rom[23983] = 8'h0b ;
            rom[23984] = 8'hf2 ;
            rom[23985] = 8'h0e ;
            rom[23986] = 8'he6 ;
            rom[23987] = 8'h14 ;
            rom[23988] = 8'h03 ;
            rom[23989] = 8'hff ;
            rom[23990] = 8'h0b ;
            rom[23991] = 8'he8 ;
            rom[23992] = 8'h00 ;
            rom[23993] = 8'hf8 ;
            rom[23994] = 8'h0a ;
            rom[23995] = 8'hf0 ;
            rom[23996] = 8'hf2 ;
            rom[23997] = 8'hdc ;
            rom[23998] = 8'hf6 ;
            rom[23999] = 8'hf9 ;
            rom[24000] = 8'hec ;
            rom[24001] = 8'h0a ;
            rom[24002] = 8'heb ;
            rom[24003] = 8'h0f ;
            rom[24004] = 8'heb ;
            rom[24005] = 8'h06 ;
            rom[24006] = 8'hdf ;
            rom[24007] = 8'hf9 ;
            rom[24008] = 8'h28 ;
            rom[24009] = 8'hf2 ;
            rom[24010] = 8'hed ;
            rom[24011] = 8'he2 ;
            rom[24012] = 8'hee ;
            rom[24013] = 8'hc4 ;
            rom[24014] = 8'he5 ;
            rom[24015] = 8'h15 ;
            rom[24016] = 8'hd5 ;
            rom[24017] = 8'he6 ;
            rom[24018] = 8'h0a ;
            rom[24019] = 8'hed ;
            rom[24020] = 8'he3 ;
            rom[24021] = 8'h05 ;
            rom[24022] = 8'hf8 ;
            rom[24023] = 8'h0c ;
            rom[24024] = 8'h05 ;
            rom[24025] = 8'hf5 ;
            rom[24026] = 8'h16 ;
            rom[24027] = 8'h18 ;
            rom[24028] = 8'h0d ;
            rom[24029] = 8'h06 ;
            rom[24030] = 8'hf6 ;
            rom[24031] = 8'he8 ;
            rom[24032] = 8'h17 ;
            rom[24033] = 8'hfb ;
            rom[24034] = 8'h08 ;
            rom[24035] = 8'he3 ;
            rom[24036] = 8'hf1 ;
            rom[24037] = 8'h11 ;
            rom[24038] = 8'he7 ;
            rom[24039] = 8'hf3 ;
            rom[24040] = 8'h03 ;
            rom[24041] = 8'h02 ;
            rom[24042] = 8'h14 ;
            rom[24043] = 8'h0d ;
            rom[24044] = 8'h25 ;
            rom[24045] = 8'hf1 ;
            rom[24046] = 8'hea ;
            rom[24047] = 8'h1d ;
            rom[24048] = 8'hf9 ;
            rom[24049] = 8'hec ;
            rom[24050] = 8'hf6 ;
            rom[24051] = 8'h1f ;
            rom[24052] = 8'hfd ;
            rom[24053] = 8'he9 ;
            rom[24054] = 8'hf7 ;
            rom[24055] = 8'hd7 ;
            rom[24056] = 8'he6 ;
            rom[24057] = 8'h17 ;
            rom[24058] = 8'hd2 ;
            rom[24059] = 8'hda ;
            rom[24060] = 8'hf7 ;
            rom[24061] = 8'h0e ;
            rom[24062] = 8'h20 ;
            rom[24063] = 8'h04 ;
            rom[24064] = 8'h0f ;
            rom[24065] = 8'he5 ;
            rom[24066] = 8'he6 ;
            rom[24067] = 8'hff ;
            rom[24068] = 8'he5 ;
            rom[24069] = 8'hdb ;
            rom[24070] = 8'h09 ;
            rom[24071] = 8'hc5 ;
            rom[24072] = 8'h28 ;
            rom[24073] = 8'h29 ;
            rom[24074] = 8'h08 ;
            rom[24075] = 8'hdc ;
            rom[24076] = 8'hf4 ;
            rom[24077] = 8'hd9 ;
            rom[24078] = 8'h0b ;
            rom[24079] = 8'hee ;
            rom[24080] = 8'h0c ;
            rom[24081] = 8'he9 ;
            rom[24082] = 8'hf2 ;
            rom[24083] = 8'h26 ;
            rom[24084] = 8'h19 ;
            rom[24085] = 8'h00 ;
            rom[24086] = 8'hcd ;
            rom[24087] = 8'hfd ;
            rom[24088] = 8'hfb ;
            rom[24089] = 8'h07 ;
            rom[24090] = 8'hfc ;
            rom[24091] = 8'hfe ;
            rom[24092] = 8'hed ;
            rom[24093] = 8'h06 ;
            rom[24094] = 8'hfb ;
            rom[24095] = 8'h17 ;
            rom[24096] = 8'hf5 ;
            rom[24097] = 8'hfc ;
            rom[24098] = 8'h0d ;
            rom[24099] = 8'hf1 ;
            rom[24100] = 8'hbd ;
            rom[24101] = 8'h00 ;
            rom[24102] = 8'hc2 ;
            rom[24103] = 8'he8 ;
            rom[24104] = 8'hcf ;
            rom[24105] = 8'he1 ;
            rom[24106] = 8'hf2 ;
            rom[24107] = 8'hf3 ;
            rom[24108] = 8'h24 ;
            rom[24109] = 8'h0b ;
            rom[24110] = 8'hde ;
            rom[24111] = 8'h0b ;
            rom[24112] = 8'hfa ;
            rom[24113] = 8'hf2 ;
            rom[24114] = 8'hf2 ;
            rom[24115] = 8'hce ;
            rom[24116] = 8'h28 ;
            rom[24117] = 8'h09 ;
            rom[24118] = 8'heb ;
            rom[24119] = 8'hf8 ;
            rom[24120] = 8'hff ;
            rom[24121] = 8'h05 ;
            rom[24122] = 8'h04 ;
            rom[24123] = 8'hea ;
            rom[24124] = 8'hf4 ;
            rom[24125] = 8'heb ;
            rom[24126] = 8'hfa ;
            rom[24127] = 8'hef ;
            rom[24128] = 8'hf0 ;
            rom[24129] = 8'h08 ;
            rom[24130] = 8'h02 ;
            rom[24131] = 8'h07 ;
            rom[24132] = 8'h22 ;
            rom[24133] = 8'h0d ;
            rom[24134] = 8'hfd ;
            rom[24135] = 8'hea ;
            rom[24136] = 8'h19 ;
            rom[24137] = 8'hd3 ;
            rom[24138] = 8'h00 ;
            rom[24139] = 8'h24 ;
            rom[24140] = 8'h28 ;
            rom[24141] = 8'hdb ;
            rom[24142] = 8'h1b ;
            rom[24143] = 8'h04 ;
            rom[24144] = 8'he9 ;
            rom[24145] = 8'hdc ;
            rom[24146] = 8'h04 ;
            rom[24147] = 8'he3 ;
            rom[24148] = 8'he4 ;
            rom[24149] = 8'hed ;
            rom[24150] = 8'hda ;
            rom[24151] = 8'h21 ;
            rom[24152] = 8'h07 ;
            rom[24153] = 8'hf6 ;
            rom[24154] = 8'h29 ;
            rom[24155] = 8'hf1 ;
            rom[24156] = 8'h03 ;
            rom[24157] = 8'h01 ;
            rom[24158] = 8'hfe ;
            rom[24159] = 8'h03 ;
            rom[24160] = 8'hd7 ;
            rom[24161] = 8'hfc ;
            rom[24162] = 8'h0a ;
            rom[24163] = 8'h2c ;
            rom[24164] = 8'hdd ;
            rom[24165] = 8'h11 ;
            rom[24166] = 8'h04 ;
            rom[24167] = 8'he5 ;
            rom[24168] = 8'h10 ;
            rom[24169] = 8'h0c ;
            rom[24170] = 8'h0b ;
            rom[24171] = 8'h11 ;
            rom[24172] = 8'h1c ;
            rom[24173] = 8'h2f ;
            rom[24174] = 8'hec ;
            rom[24175] = 8'hfb ;
            rom[24176] = 8'hee ;
            rom[24177] = 8'hec ;
            rom[24178] = 8'he9 ;
            rom[24179] = 8'he8 ;
            rom[24180] = 8'h26 ;
            rom[24181] = 8'hc8 ;
            rom[24182] = 8'h14 ;
            rom[24183] = 8'h26 ;
            rom[24184] = 8'he4 ;
            rom[24185] = 8'hfd ;
            rom[24186] = 8'he6 ;
            rom[24187] = 8'h0c ;
            rom[24188] = 8'hda ;
            rom[24189] = 8'h0a ;
            rom[24190] = 8'hd3 ;
            rom[24191] = 8'hf2 ;
            rom[24192] = 8'hf9 ;
            rom[24193] = 8'h19 ;
            rom[24194] = 8'h0d ;
            rom[24195] = 8'hc9 ;
            rom[24196] = 8'hfe ;
            rom[24197] = 8'hd4 ;
            rom[24198] = 8'hd6 ;
            rom[24199] = 8'h28 ;
            rom[24200] = 8'hec ;
            rom[24201] = 8'hfc ;
            rom[24202] = 8'hf0 ;
            rom[24203] = 8'h02 ;
            rom[24204] = 8'hcd ;
            rom[24205] = 8'h25 ;
            rom[24206] = 8'hca ;
            rom[24207] = 8'h1e ;
            rom[24208] = 8'h20 ;
            rom[24209] = 8'h05 ;
            rom[24210] = 8'h02 ;
            rom[24211] = 8'he6 ;
            rom[24212] = 8'hf9 ;
            rom[24213] = 8'hfd ;
            rom[24214] = 8'h23 ;
            rom[24215] = 8'h0b ;
            rom[24216] = 8'h12 ;
            rom[24217] = 8'h19 ;
            rom[24218] = 8'hfc ;
            rom[24219] = 8'he9 ;
            rom[24220] = 8'he4 ;
            rom[24221] = 8'h2e ;
            rom[24222] = 8'h2a ;
            rom[24223] = 8'h0e ;
            rom[24224] = 8'h21 ;
            rom[24225] = 8'he5 ;
            rom[24226] = 8'hf5 ;
            rom[24227] = 8'hd2 ;
            rom[24228] = 8'hed ;
            rom[24229] = 8'he3 ;
            rom[24230] = 8'h12 ;
            rom[24231] = 8'he4 ;
            rom[24232] = 8'hee ;
            rom[24233] = 8'hca ;
            rom[24234] = 8'he0 ;
            rom[24235] = 8'hfb ;
            rom[24236] = 8'hf3 ;
            rom[24237] = 8'hbf ;
            rom[24238] = 8'h06 ;
            rom[24239] = 8'he3 ;
            rom[24240] = 8'h0b ;
            rom[24241] = 8'hf4 ;
            rom[24242] = 8'h13 ;
            rom[24243] = 8'hf3 ;
            rom[24244] = 8'he7 ;
            rom[24245] = 8'hfa ;
            rom[24246] = 8'h0d ;
            rom[24247] = 8'heb ;
            rom[24248] = 8'hf4 ;
            rom[24249] = 8'hef ;
            rom[24250] = 8'he0 ;
            rom[24251] = 8'he2 ;
            rom[24252] = 8'h0b ;
            rom[24253] = 8'hfa ;
            rom[24254] = 8'h06 ;
            rom[24255] = 8'h0f ;
            rom[24256] = 8'h10 ;
            rom[24257] = 8'h15 ;
            rom[24258] = 8'hf5 ;
            rom[24259] = 8'hf9 ;
            rom[24260] = 8'hf2 ;
            rom[24261] = 8'hf3 ;
            rom[24262] = 8'hdc ;
            rom[24263] = 8'hec ;
            rom[24264] = 8'hd3 ;
            rom[24265] = 8'h14 ;
            rom[24266] = 8'hde ;
            rom[24267] = 8'hf2 ;
            rom[24268] = 8'hd6 ;
            rom[24269] = 8'hf1 ;
            rom[24270] = 8'hfc ;
            rom[24271] = 8'h1f ;
            rom[24272] = 8'hf2 ;
            rom[24273] = 8'h04 ;
            rom[24274] = 8'hff ;
            rom[24275] = 8'h02 ;
            rom[24276] = 8'hfe ;
            rom[24277] = 8'h02 ;
            rom[24278] = 8'he3 ;
            rom[24279] = 8'h11 ;
            rom[24280] = 8'h01 ;
            rom[24281] = 8'hf2 ;
            rom[24282] = 8'hf6 ;
            rom[24283] = 8'he2 ;
            rom[24284] = 8'h07 ;
            rom[24285] = 8'h1b ;
            rom[24286] = 8'hd2 ;
            rom[24287] = 8'hf9 ;
            rom[24288] = 8'h04 ;
            rom[24289] = 8'h1b ;
            rom[24290] = 8'hea ;
            rom[24291] = 8'hf6 ;
            rom[24292] = 8'h0b ;
            rom[24293] = 8'h12 ;
            rom[24294] = 8'h09 ;
            rom[24295] = 8'h07 ;
            rom[24296] = 8'h0c ;
            rom[24297] = 8'hfb ;
            rom[24298] = 8'he0 ;
            rom[24299] = 8'h06 ;
            rom[24300] = 8'hd3 ;
            rom[24301] = 8'hf2 ;
            rom[24302] = 8'h05 ;
            rom[24303] = 8'hf1 ;
            rom[24304] = 8'hec ;
            rom[24305] = 8'hf3 ;
            rom[24306] = 8'he5 ;
            rom[24307] = 8'h2a ;
            rom[24308] = 8'hef ;
            rom[24309] = 8'hf9 ;
            rom[24310] = 8'he8 ;
            rom[24311] = 8'hcf ;
            rom[24312] = 8'hf9 ;
            rom[24313] = 8'h1d ;
            rom[24314] = 8'hb8 ;
            rom[24315] = 8'h1b ;
            rom[24316] = 8'h03 ;
            rom[24317] = 8'hf6 ;
            rom[24318] = 8'h05 ;
            rom[24319] = 8'h3c ;
            rom[24320] = 8'hfa ;
            rom[24321] = 8'hf3 ;
            rom[24322] = 8'hfa ;
            rom[24323] = 8'he3 ;
            rom[24324] = 8'hf1 ;
            rom[24325] = 8'hf5 ;
            rom[24326] = 8'h27 ;
            rom[24327] = 8'h06 ;
            rom[24328] = 8'hed ;
            rom[24329] = 8'hf5 ;
            rom[24330] = 8'h1d ;
            rom[24331] = 8'he1 ;
            rom[24332] = 8'he8 ;
            rom[24333] = 8'hf8 ;
            rom[24334] = 8'h0f ;
            rom[24335] = 8'h01 ;
            rom[24336] = 8'h0c ;
            rom[24337] = 8'hfc ;
            rom[24338] = 8'hf3 ;
            rom[24339] = 8'h08 ;
            rom[24340] = 8'h1a ;
            rom[24341] = 8'hf1 ;
            rom[24342] = 8'hc7 ;
            rom[24343] = 8'h03 ;
            rom[24344] = 8'hd3 ;
            rom[24345] = 8'h0e ;
            rom[24346] = 8'h1c ;
            rom[24347] = 8'hf7 ;
            rom[24348] = 8'hdf ;
            rom[24349] = 8'h00 ;
            rom[24350] = 8'hf7 ;
            rom[24351] = 8'hfe ;
            rom[24352] = 8'h34 ;
            rom[24353] = 8'h0a ;
            rom[24354] = 8'hf4 ;
            rom[24355] = 8'hff ;
            rom[24356] = 8'hf2 ;
            rom[24357] = 8'h18 ;
            rom[24358] = 8'hf5 ;
            rom[24359] = 8'hed ;
            rom[24360] = 8'hf8 ;
            rom[24361] = 8'h0c ;
            rom[24362] = 8'h12 ;
            rom[24363] = 8'h0d ;
            rom[24364] = 8'h1b ;
            rom[24365] = 8'hfe ;
            rom[24366] = 8'hf7 ;
            rom[24367] = 8'hf3 ;
            rom[24368] = 8'hf6 ;
            rom[24369] = 8'hdc ;
            rom[24370] = 8'hf1 ;
            rom[24371] = 8'hc9 ;
            rom[24372] = 8'hee ;
            rom[24373] = 8'h2f ;
            rom[24374] = 8'hd3 ;
            rom[24375] = 8'h14 ;
            rom[24376] = 8'heb ;
            rom[24377] = 8'hee ;
            rom[24378] = 8'h0e ;
            rom[24379] = 8'hef ;
            rom[24380] = 8'h18 ;
            rom[24381] = 8'hed ;
            rom[24382] = 8'h1d ;
            rom[24383] = 8'hd4 ;
            rom[24384] = 8'hb9 ;
            rom[24385] = 8'h0a ;
            rom[24386] = 8'hea ;
            rom[24387] = 8'h0a ;
            rom[24388] = 8'he6 ;
            rom[24389] = 8'h20 ;
            rom[24390] = 8'hfe ;
            rom[24391] = 8'hde ;
            rom[24392] = 8'h13 ;
            rom[24393] = 8'h20 ;
            rom[24394] = 8'h0d ;
            rom[24395] = 8'h1e ;
            rom[24396] = 8'h16 ;
            rom[24397] = 8'he8 ;
            rom[24398] = 8'h1b ;
            rom[24399] = 8'h18 ;
            rom[24400] = 8'hf4 ;
            rom[24401] = 8'he1 ;
            rom[24402] = 8'h14 ;
            rom[24403] = 8'hed ;
            rom[24404] = 8'he1 ;
            rom[24405] = 8'hf2 ;
            rom[24406] = 8'hcc ;
            rom[24407] = 8'h27 ;
            rom[24408] = 8'hee ;
            rom[24409] = 8'hfb ;
            rom[24410] = 8'h09 ;
            rom[24411] = 8'h04 ;
            rom[24412] = 8'hd0 ;
            rom[24413] = 8'h02 ;
            rom[24414] = 8'h13 ;
            rom[24415] = 8'h18 ;
            rom[24416] = 8'hd6 ;
            rom[24417] = 8'heb ;
            rom[24418] = 8'hfb ;
            rom[24419] = 8'h0e ;
            rom[24420] = 8'hb7 ;
            rom[24421] = 8'h21 ;
            rom[24422] = 8'h11 ;
            rom[24423] = 8'h01 ;
            rom[24424] = 8'he1 ;
            rom[24425] = 8'h20 ;
            rom[24426] = 8'h0f ;
            rom[24427] = 8'h07 ;
            rom[24428] = 8'h18 ;
            rom[24429] = 8'he8 ;
            rom[24430] = 8'h29 ;
            rom[24431] = 8'hdd ;
            rom[24432] = 8'hfa ;
            rom[24433] = 8'hd6 ;
            rom[24434] = 8'h24 ;
            rom[24435] = 8'hff ;
            rom[24436] = 8'h1a ;
            rom[24437] = 8'h0c ;
            rom[24438] = 8'h0a ;
            rom[24439] = 8'h1d ;
            rom[24440] = 8'h11 ;
            rom[24441] = 8'hc5 ;
            rom[24442] = 8'hec ;
            rom[24443] = 8'h1c ;
            rom[24444] = 8'hb1 ;
            rom[24445] = 8'h18 ;
            rom[24446] = 8'hf5 ;
            rom[24447] = 8'hf4 ;
            rom[24448] = 8'he0 ;
            rom[24449] = 8'h09 ;
            rom[24450] = 8'h0f ;
            rom[24451] = 8'hdf ;
            rom[24452] = 8'hf7 ;
            rom[24453] = 8'hf1 ;
            rom[24454] = 8'h2c ;
            rom[24455] = 8'h08 ;
            rom[24456] = 8'h07 ;
            rom[24457] = 8'hee ;
            rom[24458] = 8'hdf ;
            rom[24459] = 8'heb ;
            rom[24460] = 8'h09 ;
            rom[24461] = 8'hf3 ;
            rom[24462] = 8'h0d ;
            rom[24463] = 8'h05 ;
            rom[24464] = 8'hb9 ;
            rom[24465] = 8'hf0 ;
            rom[24466] = 8'h19 ;
            rom[24467] = 8'h17 ;
            rom[24468] = 8'hec ;
            rom[24469] = 8'hcf ;
            rom[24470] = 8'hfb ;
            rom[24471] = 8'hd9 ;
            rom[24472] = 8'hf0 ;
            rom[24473] = 8'hec ;
            rom[24474] = 8'hcb ;
            rom[24475] = 8'h01 ;
            rom[24476] = 8'hf0 ;
            rom[24477] = 8'he9 ;
            rom[24478] = 8'hd1 ;
            rom[24479] = 8'h06 ;
            rom[24480] = 8'hd4 ;
            rom[24481] = 8'hfa ;
            rom[24482] = 8'h07 ;
            rom[24483] = 8'h16 ;
            rom[24484] = 8'h13 ;
            rom[24485] = 8'hea ;
            rom[24486] = 8'h03 ;
            rom[24487] = 8'hd6 ;
            rom[24488] = 8'h0c ;
            rom[24489] = 8'heb ;
            rom[24490] = 8'h1c ;
            rom[24491] = 8'hd7 ;
            rom[24492] = 8'hd7 ;
            rom[24493] = 8'hef ;
            rom[24494] = 8'h0c ;
            rom[24495] = 8'hc7 ;
            rom[24496] = 8'h10 ;
            rom[24497] = 8'h20 ;
            rom[24498] = 8'he2 ;
            rom[24499] = 8'he8 ;
            rom[24500] = 8'hf4 ;
            rom[24501] = 8'hfb ;
            rom[24502] = 8'hf3 ;
            rom[24503] = 8'h16 ;
            rom[24504] = 8'h11 ;
            rom[24505] = 8'h1d ;
            rom[24506] = 8'h0d ;
            rom[24507] = 8'he8 ;
            rom[24508] = 8'hf5 ;
            rom[24509] = 8'hcb ;
            rom[24510] = 8'hed ;
            rom[24511] = 8'hfa ;
            rom[24512] = 8'h28 ;
            rom[24513] = 8'h00 ;
            rom[24514] = 8'hfb ;
            rom[24515] = 8'he2 ;
            rom[24516] = 8'hf1 ;
            rom[24517] = 8'hff ;
            rom[24518] = 8'h01 ;
            rom[24519] = 8'heb ;
            rom[24520] = 8'hf8 ;
            rom[24521] = 8'hf7 ;
            rom[24522] = 8'hfa ;
            rom[24523] = 8'hf5 ;
            rom[24524] = 8'hf1 ;
            rom[24525] = 8'h11 ;
            rom[24526] = 8'hfa ;
            rom[24527] = 8'hf7 ;
            rom[24528] = 8'hf1 ;
            rom[24529] = 8'heb ;
            rom[24530] = 8'hf9 ;
            rom[24531] = 8'he4 ;
            rom[24532] = 8'h1b ;
            rom[24533] = 8'h01 ;
            rom[24534] = 8'hdf ;
            rom[24535] = 8'h01 ;
            rom[24536] = 8'he2 ;
            rom[24537] = 8'hf7 ;
            rom[24538] = 8'hd3 ;
            rom[24539] = 8'hd3 ;
            rom[24540] = 8'hcc ;
            rom[24541] = 8'he2 ;
            rom[24542] = 8'hf1 ;
            rom[24543] = 8'hf7 ;
            rom[24544] = 8'h01 ;
            rom[24545] = 8'he1 ;
            rom[24546] = 8'hf0 ;
            rom[24547] = 8'h0c ;
            rom[24548] = 8'h0f ;
            rom[24549] = 8'hd5 ;
            rom[24550] = 8'he3 ;
            rom[24551] = 8'h09 ;
            rom[24552] = 8'hed ;
            rom[24553] = 8'h0d ;
            rom[24554] = 8'haf ;
            rom[24555] = 8'hfa ;
            rom[24556] = 8'hfb ;
            rom[24557] = 8'hf1 ;
            rom[24558] = 8'h03 ;
            rom[24559] = 8'hf6 ;
            rom[24560] = 8'hf4 ;
            rom[24561] = 8'hed ;
            rom[24562] = 8'h17 ;
            rom[24563] = 8'hef ;
            rom[24564] = 8'hf5 ;
            rom[24565] = 8'hf5 ;
            rom[24566] = 8'h10 ;
            rom[24567] = 8'h02 ;
            rom[24568] = 8'hf3 ;
            rom[24569] = 8'h21 ;
            rom[24570] = 8'h02 ;
            rom[24571] = 8'h14 ;
            rom[24572] = 8'hef ;
            rom[24573] = 8'hec ;
            rom[24574] = 8'h03 ;
            rom[24575] = 8'hef ;
            rom[24576] = 8'h1b ;
            rom[24577] = 8'h01 ;
            rom[24578] = 8'h1c ;
            rom[24579] = 8'hd1 ;
            rom[24580] = 8'hfa ;
            rom[24581] = 8'h0c ;
            rom[24582] = 8'h2e ;
            rom[24583] = 8'h2f ;
            rom[24584] = 8'h04 ;
            rom[24585] = 8'h0b ;
            rom[24586] = 8'h08 ;
            rom[24587] = 8'hec ;
            rom[24588] = 8'h24 ;
            rom[24589] = 8'h13 ;
            rom[24590] = 8'h12 ;
            rom[24591] = 8'hc4 ;
            rom[24592] = 8'h14 ;
            rom[24593] = 8'he5 ;
            rom[24594] = 8'h28 ;
            rom[24595] = 8'hc9 ;
            rom[24596] = 8'h07 ;
            rom[24597] = 8'hdd ;
            rom[24598] = 8'hf6 ;
            rom[24599] = 8'hdb ;
            rom[24600] = 8'he3 ;
            rom[24601] = 8'h05 ;
            rom[24602] = 8'hee ;
            rom[24603] = 8'he0 ;
            rom[24604] = 8'hf6 ;
            rom[24605] = 8'heb ;
            rom[24606] = 8'he7 ;
            rom[24607] = 8'hdb ;
            rom[24608] = 8'hee ;
            rom[24609] = 8'h03 ;
            rom[24610] = 8'h0f ;
            rom[24611] = 8'h0c ;
            rom[24612] = 8'h1b ;
            rom[24613] = 8'h00 ;
            rom[24614] = 8'h08 ;
            rom[24615] = 8'he5 ;
            rom[24616] = 8'h05 ;
            rom[24617] = 8'he4 ;
            rom[24618] = 8'h03 ;
            rom[24619] = 8'he4 ;
            rom[24620] = 8'hf7 ;
            rom[24621] = 8'h06 ;
            rom[24622] = 8'hf5 ;
            rom[24623] = 8'hff ;
            rom[24624] = 8'h02 ;
            rom[24625] = 8'h1c ;
            rom[24626] = 8'h09 ;
            rom[24627] = 8'he5 ;
            rom[24628] = 8'hf2 ;
            rom[24629] = 8'hed ;
            rom[24630] = 8'h0b ;
            rom[24631] = 8'h01 ;
            rom[24632] = 8'hfe ;
            rom[24633] = 8'h19 ;
            rom[24634] = 8'hee ;
            rom[24635] = 8'hf0 ;
            rom[24636] = 8'he8 ;
            rom[24637] = 8'hfd ;
            rom[24638] = 8'hc9 ;
            rom[24639] = 8'hed ;
            rom[24640] = 8'h07 ;
            rom[24641] = 8'h02 ;
            rom[24642] = 8'h0d ;
            rom[24643] = 8'h07 ;
            rom[24644] = 8'hcb ;
            rom[24645] = 8'he4 ;
            rom[24646] = 8'h00 ;
            rom[24647] = 8'hf6 ;
            rom[24648] = 8'h00 ;
            rom[24649] = 8'h03 ;
            rom[24650] = 8'hf4 ;
            rom[24651] = 8'h11 ;
            rom[24652] = 8'hdc ;
            rom[24653] = 8'h04 ;
            rom[24654] = 8'h0d ;
            rom[24655] = 8'h19 ;
            rom[24656] = 8'h0a ;
            rom[24657] = 8'hfb ;
            rom[24658] = 8'hf8 ;
            rom[24659] = 8'h00 ;
            rom[24660] = 8'h08 ;
            rom[24661] = 8'h19 ;
            rom[24662] = 8'h09 ;
            rom[24663] = 8'hd9 ;
            rom[24664] = 8'hec ;
            rom[24665] = 8'hea ;
            rom[24666] = 8'hec ;
            rom[24667] = 8'hff ;
            rom[24668] = 8'hf5 ;
            rom[24669] = 8'h19 ;
            rom[24670] = 8'hd5 ;
            rom[24671] = 8'he1 ;
            rom[24672] = 8'h09 ;
            rom[24673] = 8'hfc ;
            rom[24674] = 8'h16 ;
            rom[24675] = 8'hf1 ;
            rom[24676] = 8'h00 ;
            rom[24677] = 8'he9 ;
            rom[24678] = 8'hc8 ;
            rom[24679] = 8'hfa ;
            rom[24680] = 8'h08 ;
            rom[24681] = 8'hdd ;
            rom[24682] = 8'h08 ;
            rom[24683] = 8'hfa ;
            rom[24684] = 8'h09 ;
            rom[24685] = 8'h0e ;
            rom[24686] = 8'hf7 ;
            rom[24687] = 8'hd2 ;
            rom[24688] = 8'he6 ;
            rom[24689] = 8'hb9 ;
            rom[24690] = 8'hf0 ;
            rom[24691] = 8'hfb ;
            rom[24692] = 8'h2b ;
            rom[24693] = 8'hc3 ;
            rom[24694] = 8'hec ;
            rom[24695] = 8'hef ;
            rom[24696] = 8'hf5 ;
            rom[24697] = 8'hd6 ;
            rom[24698] = 8'hf5 ;
            rom[24699] = 8'hea ;
            rom[24700] = 8'hf9 ;
            rom[24701] = 8'hf3 ;
            rom[24702] = 8'hdd ;
            rom[24703] = 8'h08 ;
            rom[24704] = 8'hf3 ;
            rom[24705] = 8'h0b ;
            rom[24706] = 8'he2 ;
            rom[24707] = 8'h06 ;
            rom[24708] = 8'hef ;
            rom[24709] = 8'hff ;
            rom[24710] = 8'he0 ;
            rom[24711] = 8'hea ;
            rom[24712] = 8'h32 ;
            rom[24713] = 8'hd4 ;
            rom[24714] = 8'h0b ;
            rom[24715] = 8'hee ;
            rom[24716] = 8'hd3 ;
            rom[24717] = 8'h0a ;
            rom[24718] = 8'h08 ;
            rom[24719] = 8'h08 ;
            rom[24720] = 8'hf8 ;
            rom[24721] = 8'hd8 ;
            rom[24722] = 8'hf6 ;
            rom[24723] = 8'hf2 ;
            rom[24724] = 8'hd5 ;
            rom[24725] = 8'heb ;
            rom[24726] = 8'hed ;
            rom[24727] = 8'hdd ;
            rom[24728] = 8'hf8 ;
            rom[24729] = 8'h11 ;
            rom[24730] = 8'hfd ;
            rom[24731] = 8'hcf ;
            rom[24732] = 8'hd9 ;
            rom[24733] = 8'hf5 ;
            rom[24734] = 8'hff ;
            rom[24735] = 8'hf6 ;
            rom[24736] = 8'hec ;
            rom[24737] = 8'hf4 ;
            rom[24738] = 8'h01 ;
            rom[24739] = 8'hfe ;
            rom[24740] = 8'hf8 ;
            rom[24741] = 8'hed ;
            rom[24742] = 8'hf8 ;
            rom[24743] = 8'hea ;
            rom[24744] = 8'h21 ;
            rom[24745] = 8'h0b ;
            rom[24746] = 8'h0a ;
            rom[24747] = 8'he8 ;
            rom[24748] = 8'he9 ;
            rom[24749] = 8'h08 ;
            rom[24750] = 8'h19 ;
            rom[24751] = 8'h02 ;
            rom[24752] = 8'hd8 ;
            rom[24753] = 8'h05 ;
            rom[24754] = 8'hde ;
            rom[24755] = 8'he6 ;
            rom[24756] = 8'hfd ;
            rom[24757] = 8'hce ;
            rom[24758] = 8'hd6 ;
            rom[24759] = 8'h03 ;
            rom[24760] = 8'h11 ;
            rom[24761] = 8'hdd ;
            rom[24762] = 8'hf1 ;
            rom[24763] = 8'hbd ;
            rom[24764] = 8'hfc ;
            rom[24765] = 8'hee ;
            rom[24766] = 8'hd1 ;
            rom[24767] = 8'h02 ;
            rom[24768] = 8'hf3 ;
            rom[24769] = 8'hee ;
            rom[24770] = 8'h0d ;
            rom[24771] = 8'hfd ;
            rom[24772] = 8'hf9 ;
            rom[24773] = 8'h16 ;
            rom[24774] = 8'h06 ;
            rom[24775] = 8'h0c ;
            rom[24776] = 8'hee ;
            rom[24777] = 8'h1a ;
            rom[24778] = 8'h07 ;
            rom[24779] = 8'hc5 ;
            rom[24780] = 8'h0d ;
            rom[24781] = 8'h11 ;
            rom[24782] = 8'h1b ;
            rom[24783] = 8'h05 ;
            rom[24784] = 8'hd1 ;
            rom[24785] = 8'hff ;
            rom[24786] = 8'hc0 ;
            rom[24787] = 8'h07 ;
            rom[24788] = 8'hea ;
            rom[24789] = 8'hcc ;
            rom[24790] = 8'hfa ;
            rom[24791] = 8'h1d ;
            rom[24792] = 8'hf1 ;
            rom[24793] = 8'he0 ;
            rom[24794] = 8'hd0 ;
            rom[24795] = 8'hdc ;
            rom[24796] = 8'hc1 ;
            rom[24797] = 8'h0e ;
            rom[24798] = 8'hf8 ;
            rom[24799] = 8'hfe ;
            rom[24800] = 8'hec ;
            rom[24801] = 8'hd6 ;
            rom[24802] = 8'hc9 ;
            rom[24803] = 8'heb ;
            rom[24804] = 8'hfb ;
            rom[24805] = 8'hf9 ;
            rom[24806] = 8'h1c ;
            rom[24807] = 8'h17 ;
            rom[24808] = 8'hd9 ;
            rom[24809] = 8'heb ;
            rom[24810] = 8'hfa ;
            rom[24811] = 8'hd4 ;
            rom[24812] = 8'h08 ;
            rom[24813] = 8'hd7 ;
            rom[24814] = 8'h01 ;
            rom[24815] = 8'h02 ;
            rom[24816] = 8'hff ;
            rom[24817] = 8'hd7 ;
            rom[24818] = 8'h20 ;
            rom[24819] = 8'h0a ;
            rom[24820] = 8'hf1 ;
            rom[24821] = 8'hf5 ;
            rom[24822] = 8'hd5 ;
            rom[24823] = 8'hbe ;
            rom[24824] = 8'hd7 ;
            rom[24825] = 8'hf3 ;
            rom[24826] = 8'h11 ;
            rom[24827] = 8'he7 ;
            rom[24828] = 8'hfd ;
            rom[24829] = 8'hd7 ;
            rom[24830] = 8'hdc ;
            rom[24831] = 8'hf1 ;
            rom[24832] = 8'h0a ;
            rom[24833] = 8'he9 ;
            rom[24834] = 8'hf3 ;
            rom[24835] = 8'h1d ;
            rom[24836] = 8'hf5 ;
            rom[24837] = 8'hdf ;
            rom[24838] = 8'h01 ;
            rom[24839] = 8'hdc ;
            rom[24840] = 8'hd6 ;
            rom[24841] = 8'hfa ;
            rom[24842] = 8'h02 ;
            rom[24843] = 8'h0d ;
            rom[24844] = 8'hf0 ;
            rom[24845] = 8'h01 ;
            rom[24846] = 8'h26 ;
            rom[24847] = 8'h0b ;
            rom[24848] = 8'h06 ;
            rom[24849] = 8'h0b ;
            rom[24850] = 8'he7 ;
            rom[24851] = 8'hf2 ;
            rom[24852] = 8'h0f ;
            rom[24853] = 8'h02 ;
            rom[24854] = 8'hd7 ;
            rom[24855] = 8'h09 ;
            rom[24856] = 8'h09 ;
            rom[24857] = 8'hf6 ;
            rom[24858] = 8'hff ;
            rom[24859] = 8'h09 ;
            rom[24860] = 8'he7 ;
            rom[24861] = 8'hec ;
            rom[24862] = 8'hd8 ;
            rom[24863] = 8'h13 ;
            rom[24864] = 8'hcb ;
            rom[24865] = 8'h21 ;
            rom[24866] = 8'hcc ;
            rom[24867] = 8'h00 ;
            rom[24868] = 8'h0b ;
            rom[24869] = 8'hd9 ;
            rom[24870] = 8'hfd ;
            rom[24871] = 8'he1 ;
            rom[24872] = 8'hb1 ;
            rom[24873] = 8'heb ;
            rom[24874] = 8'he9 ;
            rom[24875] = 8'hea ;
            rom[24876] = 8'h0a ;
            rom[24877] = 8'hf0 ;
            rom[24878] = 8'h05 ;
            rom[24879] = 8'hcb ;
            rom[24880] = 8'h18 ;
            rom[24881] = 8'hf4 ;
            rom[24882] = 8'hd6 ;
            rom[24883] = 8'heb ;
            rom[24884] = 8'h28 ;
            rom[24885] = 8'he9 ;
            rom[24886] = 8'heb ;
            rom[24887] = 8'hec ;
            rom[24888] = 8'h1b ;
            rom[24889] = 8'h00 ;
            rom[24890] = 8'hee ;
            rom[24891] = 8'h08 ;
            rom[24892] = 8'h1b ;
            rom[24893] = 8'hb9 ;
            rom[24894] = 8'hf3 ;
            rom[24895] = 8'hf7 ;
            rom[24896] = 8'hd8 ;
            rom[24897] = 8'h15 ;
            rom[24898] = 8'h14 ;
            rom[24899] = 8'h10 ;
            rom[24900] = 8'hc7 ;
            rom[24901] = 8'heb ;
            rom[24902] = 8'he6 ;
            rom[24903] = 8'hfa ;
            rom[24904] = 8'hfc ;
            rom[24905] = 8'hfa ;
            rom[24906] = 8'h06 ;
            rom[24907] = 8'h1b ;
            rom[24908] = 8'h0f ;
            rom[24909] = 8'h1d ;
            rom[24910] = 8'hc1 ;
            rom[24911] = 8'h16 ;
            rom[24912] = 8'he7 ;
            rom[24913] = 8'he9 ;
            rom[24914] = 8'hec ;
            rom[24915] = 8'hfe ;
            rom[24916] = 8'hf7 ;
            rom[24917] = 8'hfe ;
            rom[24918] = 8'hef ;
            rom[24919] = 8'h08 ;
            rom[24920] = 8'h07 ;
            rom[24921] = 8'he6 ;
            rom[24922] = 8'hfa ;
            rom[24923] = 8'h11 ;
            rom[24924] = 8'h13 ;
            rom[24925] = 8'h04 ;
            rom[24926] = 8'h03 ;
            rom[24927] = 8'h03 ;
            rom[24928] = 8'h09 ;
            rom[24929] = 8'hd4 ;
            rom[24930] = 8'h12 ;
            rom[24931] = 8'heb ;
            rom[24932] = 8'he0 ;
            rom[24933] = 8'hd0 ;
            rom[24934] = 8'h14 ;
            rom[24935] = 8'h12 ;
            rom[24936] = 8'hcd ;
            rom[24937] = 8'hd3 ;
            rom[24938] = 8'hf9 ;
            rom[24939] = 8'hef ;
            rom[24940] = 8'hef ;
            rom[24941] = 8'he3 ;
            rom[24942] = 8'h19 ;
            rom[24943] = 8'h21 ;
            rom[24944] = 8'h25 ;
            rom[24945] = 8'h10 ;
            rom[24946] = 8'h08 ;
            rom[24947] = 8'h10 ;
            rom[24948] = 8'hf8 ;
            rom[24949] = 8'hfe ;
            rom[24950] = 8'h1b ;
            rom[24951] = 8'h0d ;
            rom[24952] = 8'he9 ;
            rom[24953] = 8'h08 ;
            rom[24954] = 8'hfa ;
            rom[24955] = 8'hc5 ;
            rom[24956] = 8'hfd ;
            rom[24957] = 8'h07 ;
            rom[24958] = 8'hc0 ;
            rom[24959] = 8'hd3 ;
            rom[24960] = 8'hf7 ;
            rom[24961] = 8'hfe ;
            rom[24962] = 8'h0a ;
            rom[24963] = 8'h0b ;
            rom[24964] = 8'hcf ;
            rom[24965] = 8'hf5 ;
            rom[24966] = 8'h0f ;
            rom[24967] = 8'hdc ;
            rom[24968] = 8'hea ;
            rom[24969] = 8'h18 ;
            rom[24970] = 8'hc3 ;
            rom[24971] = 8'h06 ;
            rom[24972] = 8'h0e ;
            rom[24973] = 8'hed ;
            rom[24974] = 8'hde ;
            rom[24975] = 8'h17 ;
            rom[24976] = 8'h29 ;
            rom[24977] = 8'he7 ;
            rom[24978] = 8'h1d ;
            rom[24979] = 8'h0e ;
            rom[24980] = 8'hff ;
            rom[24981] = 8'hdc ;
            rom[24982] = 8'hd5 ;
            rom[24983] = 8'h2f ;
            rom[24984] = 8'hfc ;
            rom[24985] = 8'h0f ;
            rom[24986] = 8'hf1 ;
            rom[24987] = 8'hfb ;
            rom[24988] = 8'hd8 ;
            rom[24989] = 8'h13 ;
            rom[24990] = 8'h0c ;
            rom[24991] = 8'hd8 ;
            rom[24992] = 8'hf3 ;
            rom[24993] = 8'hf9 ;
            rom[24994] = 8'h0b ;
            rom[24995] = 8'hd4 ;
            rom[24996] = 8'hf7 ;
            rom[24997] = 8'hef ;
            rom[24998] = 8'h16 ;
            rom[24999] = 8'h0f ;
            rom[25000] = 8'hf3 ;
            rom[25001] = 8'hdc ;
            rom[25002] = 8'h02 ;
            rom[25003] = 8'hfe ;
            rom[25004] = 8'hf0 ;
            rom[25005] = 8'he9 ;
            rom[25006] = 8'h07 ;
            rom[25007] = 8'hce ;
            rom[25008] = 8'h05 ;
            rom[25009] = 8'hf3 ;
            rom[25010] = 8'hfc ;
            rom[25011] = 8'h1f ;
            rom[25012] = 8'hf1 ;
            rom[25013] = 8'hf8 ;
            rom[25014] = 8'h08 ;
            rom[25015] = 8'hc9 ;
            rom[25016] = 8'h09 ;
            rom[25017] = 8'h1c ;
            rom[25018] = 8'h0b ;
            rom[25019] = 8'h0f ;
            rom[25020] = 8'hf0 ;
            rom[25021] = 8'h09 ;
            rom[25022] = 8'hcc ;
            rom[25023] = 8'h01 ;
            rom[25024] = 8'hfe ;
            rom[25025] = 8'he2 ;
            rom[25026] = 8'hde ;
            rom[25027] = 8'hf4 ;
            rom[25028] = 8'hdb ;
            rom[25029] = 8'hf2 ;
            rom[25030] = 8'hf0 ;
            rom[25031] = 8'hd6 ;
            rom[25032] = 8'hb8 ;
            rom[25033] = 8'hcf ;
            rom[25034] = 8'h23 ;
            rom[25035] = 8'h14 ;
            rom[25036] = 8'hf3 ;
            rom[25037] = 8'h07 ;
            rom[25038] = 8'hd1 ;
            rom[25039] = 8'h07 ;
            rom[25040] = 8'hf8 ;
            rom[25041] = 8'hd5 ;
            rom[25042] = 8'hef ;
            rom[25043] = 8'hf3 ;
            rom[25044] = 8'h05 ;
            rom[25045] = 8'h02 ;
            rom[25046] = 8'hff ;
            rom[25047] = 8'hef ;
            rom[25048] = 8'h0c ;
            rom[25049] = 8'h18 ;
            rom[25050] = 8'h08 ;
            rom[25051] = 8'h12 ;
            rom[25052] = 8'hdb ;
            rom[25053] = 8'hd8 ;
            rom[25054] = 8'hfc ;
            rom[25055] = 8'h06 ;
            rom[25056] = 8'h20 ;
            rom[25057] = 8'hf2 ;
            rom[25058] = 8'hdb ;
            rom[25059] = 8'h10 ;
            rom[25060] = 8'h2d ;
            rom[25061] = 8'hed ;
            rom[25062] = 8'h06 ;
            rom[25063] = 8'hdb ;
            rom[25064] = 8'hff ;
            rom[25065] = 8'hbc ;
            rom[25066] = 8'h02 ;
            rom[25067] = 8'h11 ;
            rom[25068] = 8'hd5 ;
            rom[25069] = 8'hf0 ;
            rom[25070] = 8'h00 ;
            rom[25071] = 8'he2 ;
            rom[25072] = 8'h0b ;
            rom[25073] = 8'hed ;
            rom[25074] = 8'h15 ;
            rom[25075] = 8'he4 ;
            rom[25076] = 8'he0 ;
            rom[25077] = 8'hce ;
            rom[25078] = 8'hef ;
            rom[25079] = 8'he8 ;
            rom[25080] = 8'hdf ;
            rom[25081] = 8'hf6 ;
            rom[25082] = 8'h01 ;
            rom[25083] = 8'h09 ;
            rom[25084] = 8'heb ;
            rom[25085] = 8'hbc ;
            rom[25086] = 8'hea ;
            rom[25087] = 8'h08 ;
            rom[25088] = 8'hf2 ;
            rom[25089] = 8'h04 ;
            rom[25090] = 8'hfa ;
            rom[25091] = 8'h0e ;
            rom[25092] = 8'h20 ;
            rom[25093] = 8'he1 ;
            rom[25094] = 8'h06 ;
            rom[25095] = 8'hfc ;
            rom[25096] = 8'h02 ;
            rom[25097] = 8'hfe ;
            rom[25098] = 8'heb ;
            rom[25099] = 8'he3 ;
            rom[25100] = 8'hd5 ;
            rom[25101] = 8'h01 ;
            rom[25102] = 8'hec ;
            rom[25103] = 8'he9 ;
            rom[25104] = 8'hcc ;
            rom[25105] = 8'h01 ;
            rom[25106] = 8'he6 ;
            rom[25107] = 8'hc2 ;
            rom[25108] = 8'h11 ;
            rom[25109] = 8'h04 ;
            rom[25110] = 8'h0e ;
            rom[25111] = 8'h11 ;
            rom[25112] = 8'h0e ;
            rom[25113] = 8'hf6 ;
            rom[25114] = 8'he9 ;
            rom[25115] = 8'h2d ;
            rom[25116] = 8'h1b ;
            rom[25117] = 8'he1 ;
            rom[25118] = 8'h3d ;
            rom[25119] = 8'h02 ;
            rom[25120] = 8'hf3 ;
            rom[25121] = 8'hed ;
            rom[25122] = 8'h0c ;
            rom[25123] = 8'hfd ;
            rom[25124] = 8'h10 ;
            rom[25125] = 8'h03 ;
            rom[25126] = 8'hfc ;
            rom[25127] = 8'h15 ;
            rom[25128] = 8'hce ;
            rom[25129] = 8'h0c ;
            rom[25130] = 8'hf9 ;
            rom[25131] = 8'h00 ;
            rom[25132] = 8'h08 ;
            rom[25133] = 8'h01 ;
            rom[25134] = 8'hb7 ;
            rom[25135] = 8'h1c ;
            rom[25136] = 8'h09 ;
            rom[25137] = 8'hfe ;
            rom[25138] = 8'hd9 ;
            rom[25139] = 8'hd8 ;
            rom[25140] = 8'hd9 ;
            rom[25141] = 8'h02 ;
            rom[25142] = 8'hcf ;
            rom[25143] = 8'h25 ;
            rom[25144] = 8'hf9 ;
            rom[25145] = 8'hf6 ;
            rom[25146] = 8'hf3 ;
            rom[25147] = 8'hfc ;
            rom[25148] = 8'h1a ;
            rom[25149] = 8'hfc ;
            rom[25150] = 8'hdf ;
            rom[25151] = 8'hf6 ;
            rom[25152] = 8'h07 ;
            rom[25153] = 8'h12 ;
            rom[25154] = 8'he3 ;
            rom[25155] = 8'h01 ;
            rom[25156] = 8'h20 ;
            rom[25157] = 8'h0b ;
            rom[25158] = 8'hf1 ;
            rom[25159] = 8'hf8 ;
            rom[25160] = 8'h16 ;
            rom[25161] = 8'h03 ;
            rom[25162] = 8'hef ;
            rom[25163] = 8'hff ;
            rom[25164] = 8'hf8 ;
            rom[25165] = 8'h0b ;
            rom[25166] = 8'hdb ;
            rom[25167] = 8'he4 ;
            rom[25168] = 8'hfe ;
            rom[25169] = 8'h12 ;
            rom[25170] = 8'he7 ;
            rom[25171] = 8'hf8 ;
            rom[25172] = 8'hf7 ;
            rom[25173] = 8'hef ;
            rom[25174] = 8'h1a ;
            rom[25175] = 8'hfd ;
            rom[25176] = 8'hf9 ;
            rom[25177] = 8'h13 ;
            rom[25178] = 8'hfe ;
            rom[25179] = 8'hc8 ;
            rom[25180] = 8'h26 ;
            rom[25181] = 8'h01 ;
            rom[25182] = 8'hdb ;
            rom[25183] = 8'hdf ;
            rom[25184] = 8'hd1 ;
            rom[25185] = 8'h09 ;
            rom[25186] = 8'hf7 ;
            rom[25187] = 8'h0b ;
            rom[25188] = 8'he2 ;
            rom[25189] = 8'h25 ;
            rom[25190] = 8'h14 ;
            rom[25191] = 8'heb ;
            rom[25192] = 8'hd6 ;
            rom[25193] = 8'h1e ;
            rom[25194] = 8'hf7 ;
            rom[25195] = 8'hdc ;
            rom[25196] = 8'hbc ;
            rom[25197] = 8'hfd ;
            rom[25198] = 8'he1 ;
            rom[25199] = 8'h0b ;
            rom[25200] = 8'he8 ;
            rom[25201] = 8'h19 ;
            rom[25202] = 8'h02 ;
            rom[25203] = 8'hed ;
            rom[25204] = 8'he3 ;
            rom[25205] = 8'hfc ;
            rom[25206] = 8'h04 ;
            rom[25207] = 8'h07 ;
            rom[25208] = 8'hf9 ;
            rom[25209] = 8'hfe ;
            rom[25210] = 8'hd2 ;
            rom[25211] = 8'h2a ;
            rom[25212] = 8'hec ;
            rom[25213] = 8'h16 ;
            rom[25214] = 8'h13 ;
            rom[25215] = 8'he4 ;
            rom[25216] = 8'hf2 ;
            rom[25217] = 8'hdf ;
            rom[25218] = 8'h05 ;
            rom[25219] = 8'he9 ;
            rom[25220] = 8'h1c ;
            rom[25221] = 8'hc8 ;
            rom[25222] = 8'hf4 ;
            rom[25223] = 8'h07 ;
            rom[25224] = 8'h02 ;
            rom[25225] = 8'hf9 ;
            rom[25226] = 8'h25 ;
            rom[25227] = 8'hc6 ;
            rom[25228] = 8'h0f ;
            rom[25229] = 8'h15 ;
            rom[25230] = 8'h10 ;
            rom[25231] = 8'hfa ;
            rom[25232] = 8'h06 ;
            rom[25233] = 8'hd3 ;
            rom[25234] = 8'h0e ;
            rom[25235] = 8'hf8 ;
            rom[25236] = 8'hfb ;
            rom[25237] = 8'h23 ;
            rom[25238] = 8'hf0 ;
            rom[25239] = 8'h14 ;
            rom[25240] = 8'h1c ;
            rom[25241] = 8'h12 ;
            rom[25242] = 8'h25 ;
            rom[25243] = 8'h03 ;
            rom[25244] = 8'hc5 ;
            rom[25245] = 8'h06 ;
            rom[25246] = 8'h09 ;
            rom[25247] = 8'hff ;
            rom[25248] = 8'h02 ;
            rom[25249] = 8'he8 ;
            rom[25250] = 8'hea ;
            rom[25251] = 8'h0e ;
            rom[25252] = 8'h07 ;
            rom[25253] = 8'hf9 ;
            rom[25254] = 8'he7 ;
            rom[25255] = 8'hfc ;
            rom[25256] = 8'h07 ;
            rom[25257] = 8'hf2 ;
            rom[25258] = 8'h0d ;
            rom[25259] = 8'hef ;
            rom[25260] = 8'hd6 ;
            rom[25261] = 8'h28 ;
            rom[25262] = 8'h10 ;
            rom[25263] = 8'hd2 ;
            rom[25264] = 8'hd1 ;
            rom[25265] = 8'h14 ;
            rom[25266] = 8'h08 ;
            rom[25267] = 8'he5 ;
            rom[25268] = 8'hea ;
            rom[25269] = 8'hf9 ;
            rom[25270] = 8'h08 ;
            rom[25271] = 8'h24 ;
            rom[25272] = 8'hfb ;
            rom[25273] = 8'h10 ;
            rom[25274] = 8'h18 ;
            rom[25275] = 8'h05 ;
            rom[25276] = 8'hdc ;
            rom[25277] = 8'he7 ;
            rom[25278] = 8'hf1 ;
            rom[25279] = 8'he3 ;
            rom[25280] = 8'h0b ;
            rom[25281] = 8'hfc ;
            rom[25282] = 8'hea ;
            rom[25283] = 8'hff ;
            rom[25284] = 8'hf7 ;
            rom[25285] = 8'h10 ;
            rom[25286] = 8'hff ;
            rom[25287] = 8'hff ;
            rom[25288] = 8'h06 ;
            rom[25289] = 8'hce ;
            rom[25290] = 8'hea ;
            rom[25291] = 8'hfd ;
            rom[25292] = 8'h0c ;
            rom[25293] = 8'hf6 ;
            rom[25294] = 8'hc0 ;
            rom[25295] = 8'h16 ;
            rom[25296] = 8'hf8 ;
            rom[25297] = 8'hd0 ;
            rom[25298] = 8'h02 ;
            rom[25299] = 8'h1d ;
            rom[25300] = 8'h0f ;
            rom[25301] = 8'h09 ;
            rom[25302] = 8'h03 ;
            rom[25303] = 8'hea ;
            rom[25304] = 8'hdf ;
            rom[25305] = 8'h08 ;
            rom[25306] = 8'h03 ;
            rom[25307] = 8'hf4 ;
            rom[25308] = 8'h00 ;
            rom[25309] = 8'h18 ;
            rom[25310] = 8'h13 ;
            rom[25311] = 8'hff ;
            rom[25312] = 8'hfa ;
            rom[25313] = 8'hfd ;
            rom[25314] = 8'h1c ;
            rom[25315] = 8'hef ;
            rom[25316] = 8'hfa ;
            rom[25317] = 8'h0c ;
            rom[25318] = 8'h1c ;
            rom[25319] = 8'hc7 ;
            rom[25320] = 8'hfe ;
            rom[25321] = 8'hd0 ;
            rom[25322] = 8'hde ;
            rom[25323] = 8'h1b ;
            rom[25324] = 8'he3 ;
            rom[25325] = 8'h08 ;
            rom[25326] = 8'h09 ;
            rom[25327] = 8'hfc ;
            rom[25328] = 8'h02 ;
            rom[25329] = 8'hfb ;
            rom[25330] = 8'h10 ;
            rom[25331] = 8'hf7 ;
            rom[25332] = 8'hf9 ;
            rom[25333] = 8'h0a ;
            rom[25334] = 8'hc4 ;
            rom[25335] = 8'he0 ;
            rom[25336] = 8'hcb ;
            rom[25337] = 8'h22 ;
            rom[25338] = 8'h18 ;
            rom[25339] = 8'h04 ;
            rom[25340] = 8'he5 ;
            rom[25341] = 8'he5 ;
            rom[25342] = 8'he4 ;
            rom[25343] = 8'hfb ;
            rom[25344] = 8'hec ;
            rom[25345] = 8'hc7 ;
            rom[25346] = 8'he4 ;
            rom[25347] = 8'h07 ;
            rom[25348] = 8'hb5 ;
            rom[25349] = 8'h0e ;
            rom[25350] = 8'h10 ;
            rom[25351] = 8'h0e ;
            rom[25352] = 8'h10 ;
            rom[25353] = 8'hcb ;
            rom[25354] = 8'heb ;
            rom[25355] = 8'hfe ;
            rom[25356] = 8'h08 ;
            rom[25357] = 8'he0 ;
            rom[25358] = 8'h0b ;
            rom[25359] = 8'hd0 ;
            rom[25360] = 8'h02 ;
            rom[25361] = 8'hfb ;
            rom[25362] = 8'he4 ;
            rom[25363] = 8'hd6 ;
            rom[25364] = 8'h04 ;
            rom[25365] = 8'hf6 ;
            rom[25366] = 8'hdf ;
            rom[25367] = 8'h08 ;
            rom[25368] = 8'h11 ;
            rom[25369] = 8'hc6 ;
            rom[25370] = 8'he6 ;
            rom[25371] = 8'h00 ;
            rom[25372] = 8'hfa ;
            rom[25373] = 8'h2f ;
            rom[25374] = 8'he4 ;
            rom[25375] = 8'h0b ;
            rom[25376] = 8'h0b ;
            rom[25377] = 8'hf3 ;
            rom[25378] = 8'hed ;
            rom[25379] = 8'h03 ;
            rom[25380] = 8'h16 ;
            rom[25381] = 8'h27 ;
            rom[25382] = 8'h16 ;
            rom[25383] = 8'hcb ;
            rom[25384] = 8'hf5 ;
            rom[25385] = 8'hfc ;
            rom[25386] = 8'h13 ;
            rom[25387] = 8'hf8 ;
            rom[25388] = 8'h19 ;
            rom[25389] = 8'hfe ;
            rom[25390] = 8'hf0 ;
            rom[25391] = 8'h18 ;
            rom[25392] = 8'hf2 ;
            rom[25393] = 8'h11 ;
            rom[25394] = 8'hff ;
            rom[25395] = 8'hee ;
            rom[25396] = 8'h26 ;
            rom[25397] = 8'h0c ;
            rom[25398] = 8'hf1 ;
            rom[25399] = 8'h03 ;
            rom[25400] = 8'hf5 ;
            rom[25401] = 8'hd8 ;
            rom[25402] = 8'hce ;
            rom[25403] = 8'hf8 ;
            rom[25404] = 8'h05 ;
            rom[25405] = 8'hff ;
            rom[25406] = 8'h12 ;
            rom[25407] = 8'hed ;
            rom[25408] = 8'h14 ;
            rom[25409] = 8'h1a ;
            rom[25410] = 8'hfa ;
            rom[25411] = 8'h09 ;
            rom[25412] = 8'hfb ;
            rom[25413] = 8'h19 ;
            rom[25414] = 8'hef ;
            rom[25415] = 8'hf3 ;
            rom[25416] = 8'hf6 ;
            rom[25417] = 8'h13 ;
            rom[25418] = 8'hea ;
            rom[25419] = 8'h0f ;
            rom[25420] = 8'hc5 ;
            rom[25421] = 8'h1c ;
            rom[25422] = 8'hf4 ;
            rom[25423] = 8'h02 ;
            rom[25424] = 8'hdd ;
            rom[25425] = 8'hfd ;
            rom[25426] = 8'h05 ;
            rom[25427] = 8'hec ;
            rom[25428] = 8'hea ;
            rom[25429] = 8'h07 ;
            rom[25430] = 8'hd1 ;
            rom[25431] = 8'h12 ;
            rom[25432] = 8'h1d ;
            rom[25433] = 8'h03 ;
            rom[25434] = 8'h05 ;
            rom[25435] = 8'h01 ;
            rom[25436] = 8'h03 ;
            rom[25437] = 8'hec ;
            rom[25438] = 8'hfe ;
            rom[25439] = 8'h03 ;
            rom[25440] = 8'hc4 ;
            rom[25441] = 8'h2f ;
            rom[25442] = 8'he3 ;
            rom[25443] = 8'h18 ;
            rom[25444] = 8'hbd ;
            rom[25445] = 8'he9 ;
            rom[25446] = 8'hf5 ;
            rom[25447] = 8'hf7 ;
            rom[25448] = 8'h04 ;
            rom[25449] = 8'h01 ;
            rom[25450] = 8'hf9 ;
            rom[25451] = 8'h10 ;
            rom[25452] = 8'h14 ;
            rom[25453] = 8'hfe ;
            rom[25454] = 8'hda ;
            rom[25455] = 8'h07 ;
            rom[25456] = 8'h00 ;
            rom[25457] = 8'h11 ;
            rom[25458] = 8'hf4 ;
            rom[25459] = 8'h24 ;
            rom[25460] = 8'h0e ;
            rom[25461] = 8'h09 ;
            rom[25462] = 8'h11 ;
            rom[25463] = 8'h0b ;
            rom[25464] = 8'hf3 ;
            rom[25465] = 8'hf9 ;
            rom[25466] = 8'he5 ;
            rom[25467] = 8'h11 ;
            rom[25468] = 8'h17 ;
            rom[25469] = 8'h1e ;
            rom[25470] = 8'h04 ;
            rom[25471] = 8'hf8 ;
            rom[25472] = 8'h21 ;
            rom[25473] = 8'hc3 ;
            rom[25474] = 8'hc8 ;
            rom[25475] = 8'h32 ;
            rom[25476] = 8'h04 ;
            rom[25477] = 8'hf3 ;
            rom[25478] = 8'h1d ;
            rom[25479] = 8'hfa ;
            rom[25480] = 8'he5 ;
            rom[25481] = 8'hfe ;
            rom[25482] = 8'hfc ;
            rom[25483] = 8'hd6 ;
            rom[25484] = 8'heb ;
            rom[25485] = 8'hd2 ;
            rom[25486] = 8'hf8 ;
            rom[25487] = 8'hd4 ;
            rom[25488] = 8'hf9 ;
            rom[25489] = 8'hd1 ;
            rom[25490] = 8'h01 ;
            rom[25491] = 8'hfe ;
            rom[25492] = 8'h07 ;
            rom[25493] = 8'hf2 ;
            rom[25494] = 8'h0e ;
            rom[25495] = 8'h17 ;
            rom[25496] = 8'h14 ;
            rom[25497] = 8'h07 ;
            rom[25498] = 8'he7 ;
            rom[25499] = 8'h20 ;
            rom[25500] = 8'h0e ;
            rom[25501] = 8'h33 ;
            rom[25502] = 8'h02 ;
            rom[25503] = 8'h05 ;
            rom[25504] = 8'h0d ;
            rom[25505] = 8'hf7 ;
            rom[25506] = 8'hf1 ;
            rom[25507] = 8'h0a ;
            rom[25508] = 8'hcd ;
            rom[25509] = 8'hfa ;
            rom[25510] = 8'h06 ;
            rom[25511] = 8'hf7 ;
            rom[25512] = 8'hff ;
            rom[25513] = 8'h15 ;
            rom[25514] = 8'h15 ;
            rom[25515] = 8'hca ;
            rom[25516] = 8'h25 ;
            rom[25517] = 8'h11 ;
            rom[25518] = 8'hb9 ;
            rom[25519] = 8'h18 ;
            rom[25520] = 8'h0d ;
            rom[25521] = 8'he7 ;
            rom[25522] = 8'h1e ;
            rom[25523] = 8'h00 ;
            rom[25524] = 8'h11 ;
            rom[25525] = 8'hf0 ;
            rom[25526] = 8'h0f ;
            rom[25527] = 8'h0b ;
            rom[25528] = 8'he9 ;
            rom[25529] = 8'h1b ;
            rom[25530] = 8'h12 ;
            rom[25531] = 8'h06 ;
            rom[25532] = 8'h0d ;
            rom[25533] = 8'h02 ;
            rom[25534] = 8'hd7 ;
            rom[25535] = 8'hdf ;
            rom[25536] = 8'h10 ;
            rom[25537] = 8'h16 ;
            rom[25538] = 8'h0f ;
            rom[25539] = 8'hf2 ;
            rom[25540] = 8'h07 ;
            rom[25541] = 8'hd7 ;
            rom[25542] = 8'hfa ;
            rom[25543] = 8'hfa ;
            rom[25544] = 8'hf0 ;
            rom[25545] = 8'hfa ;
            rom[25546] = 8'h18 ;
            rom[25547] = 8'h05 ;
            rom[25548] = 8'he2 ;
            rom[25549] = 8'hf2 ;
            rom[25550] = 8'hd9 ;
            rom[25551] = 8'hf7 ;
            rom[25552] = 8'hec ;
            rom[25553] = 8'hcc ;
            rom[25554] = 8'he7 ;
            rom[25555] = 8'hfa ;
            rom[25556] = 8'hd6 ;
            rom[25557] = 8'h01 ;
            rom[25558] = 8'h02 ;
            rom[25559] = 8'h36 ;
            rom[25560] = 8'hda ;
            rom[25561] = 8'h0c ;
            rom[25562] = 8'h09 ;
            rom[25563] = 8'h15 ;
            rom[25564] = 8'hfc ;
            rom[25565] = 8'hef ;
            rom[25566] = 8'he9 ;
            rom[25567] = 8'hfa ;
            rom[25568] = 8'h16 ;
            rom[25569] = 8'h16 ;
            rom[25570] = 8'hbf ;
            rom[25571] = 8'hea ;
            rom[25572] = 8'h09 ;
            rom[25573] = 8'hf9 ;
            rom[25574] = 8'hd3 ;
            rom[25575] = 8'hdb ;
            rom[25576] = 8'hf5 ;
            rom[25577] = 8'h09 ;
            rom[25578] = 8'h16 ;
            rom[25579] = 8'h1f ;
            rom[25580] = 8'h12 ;
            rom[25581] = 8'hfb ;
            rom[25582] = 8'hed ;
            rom[25583] = 8'h07 ;
            rom[25584] = 8'h02 ;
            rom[25585] = 8'hf0 ;
            rom[25586] = 8'h06 ;
            rom[25587] = 8'h1f ;
            rom[25588] = 8'hcc ;
            rom[25589] = 8'h12 ;
            rom[25590] = 8'h03 ;
            rom[25591] = 8'hdc ;
            rom[25592] = 8'h06 ;
            rom[25593] = 8'hf2 ;
            rom[25594] = 8'hf0 ;
            rom[25595] = 8'h0c ;
            rom[25596] = 8'h14 ;
            rom[25597] = 8'hf2 ;
            rom[25598] = 8'h1c ;
            rom[25599] = 8'h07 ;
            rom[25600] = 8'h0a ;
            rom[25601] = 8'h23 ;
            rom[25602] = 8'hf1 ;
            rom[25603] = 8'hf4 ;
            rom[25604] = 8'h04 ;
            rom[25605] = 8'he6 ;
            rom[25606] = 8'hea ;
            rom[25607] = 8'he4 ;
            rom[25608] = 8'h1f ;
            rom[25609] = 8'he2 ;
            rom[25610] = 8'hea ;
            rom[25611] = 8'hff ;
            rom[25612] = 8'he7 ;
            rom[25613] = 8'hff ;
            rom[25614] = 8'h06 ;
            rom[25615] = 8'hfd ;
            rom[25616] = 8'hc0 ;
            rom[25617] = 8'h0b ;
            rom[25618] = 8'h0a ;
            rom[25619] = 8'he9 ;
            rom[25620] = 8'hf1 ;
            rom[25621] = 8'h03 ;
            rom[25622] = 8'h05 ;
            rom[25623] = 8'hf4 ;
            rom[25624] = 8'hca ;
            rom[25625] = 8'hda ;
            rom[25626] = 8'hf8 ;
            rom[25627] = 8'hf9 ;
            rom[25628] = 8'hf7 ;
            rom[25629] = 8'h17 ;
            rom[25630] = 8'h02 ;
            rom[25631] = 8'he8 ;
            rom[25632] = 8'hf8 ;
            rom[25633] = 8'hfc ;
            rom[25634] = 8'h0f ;
            rom[25635] = 8'h11 ;
            rom[25636] = 8'hf0 ;
            rom[25637] = 8'h01 ;
            rom[25638] = 8'hf7 ;
            rom[25639] = 8'hec ;
            rom[25640] = 8'h04 ;
            rom[25641] = 8'hfe ;
            rom[25642] = 8'h3a ;
            rom[25643] = 8'h16 ;
            rom[25644] = 8'hfb ;
            rom[25645] = 8'hfc ;
            rom[25646] = 8'h0a ;
            rom[25647] = 8'hf7 ;
            rom[25648] = 8'hfa ;
            rom[25649] = 8'h0e ;
            rom[25650] = 8'hf5 ;
            rom[25651] = 8'hc8 ;
            rom[25652] = 8'hf8 ;
            rom[25653] = 8'hf0 ;
            rom[25654] = 8'hec ;
            rom[25655] = 8'h0f ;
            rom[25656] = 8'h2f ;
            rom[25657] = 8'hcf ;
            rom[25658] = 8'hea ;
            rom[25659] = 8'he5 ;
            rom[25660] = 8'h17 ;
            rom[25661] = 8'h12 ;
            rom[25662] = 8'h17 ;
            rom[25663] = 8'hb8 ;
            rom[25664] = 8'h01 ;
            rom[25665] = 8'hff ;
            rom[25666] = 8'hf1 ;
            rom[25667] = 8'hf5 ;
            rom[25668] = 8'hf5 ;
            rom[25669] = 8'h12 ;
            rom[25670] = 8'he0 ;
            rom[25671] = 8'h2a ;
            rom[25672] = 8'h09 ;
            rom[25673] = 8'h08 ;
            rom[25674] = 8'hd0 ;
            rom[25675] = 8'hd4 ;
            rom[25676] = 8'hf4 ;
            rom[25677] = 8'hfd ;
            rom[25678] = 8'he8 ;
            rom[25679] = 8'he6 ;
            rom[25680] = 8'hec ;
            rom[25681] = 8'hfe ;
            rom[25682] = 8'h07 ;
            rom[25683] = 8'h0d ;
            rom[25684] = 8'hf4 ;
            rom[25685] = 8'hf3 ;
            rom[25686] = 8'hf3 ;
            rom[25687] = 8'hf8 ;
            rom[25688] = 8'hc9 ;
            rom[25689] = 8'h11 ;
            rom[25690] = 8'he8 ;
            rom[25691] = 8'hf4 ;
            rom[25692] = 8'hf4 ;
            rom[25693] = 8'h07 ;
            rom[25694] = 8'hfa ;
            rom[25695] = 8'hfb ;
            rom[25696] = 8'he3 ;
            rom[25697] = 8'h0a ;
            rom[25698] = 8'hf5 ;
            rom[25699] = 8'h07 ;
            rom[25700] = 8'hf8 ;
            rom[25701] = 8'hf9 ;
            rom[25702] = 8'h05 ;
            rom[25703] = 8'hd0 ;
            rom[25704] = 8'hf8 ;
            rom[25705] = 8'h18 ;
            rom[25706] = 8'he4 ;
            rom[25707] = 8'hec ;
            rom[25708] = 8'h1a ;
            rom[25709] = 8'hee ;
            rom[25710] = 8'he3 ;
            rom[25711] = 8'hff ;
            rom[25712] = 8'hd8 ;
            rom[25713] = 8'h01 ;
            rom[25714] = 8'hf3 ;
            rom[25715] = 8'h23 ;
            rom[25716] = 8'hf2 ;
            rom[25717] = 8'h15 ;
            rom[25718] = 8'hed ;
            rom[25719] = 8'h0c ;
            rom[25720] = 8'hed ;
            rom[25721] = 8'hf6 ;
            rom[25722] = 8'he2 ;
            rom[25723] = 8'hfb ;
            rom[25724] = 8'hf6 ;
            rom[25725] = 8'hfb ;
            rom[25726] = 8'h0c ;
            rom[25727] = 8'he4 ;
            rom[25728] = 8'he7 ;
            rom[25729] = 8'heb ;
            rom[25730] = 8'h0c ;
            rom[25731] = 8'hbe ;
            rom[25732] = 8'h00 ;
            rom[25733] = 8'hf3 ;
            rom[25734] = 8'h1f ;
            rom[25735] = 8'h11 ;
            rom[25736] = 8'hfd ;
            rom[25737] = 8'hc9 ;
            rom[25738] = 8'h0c ;
            rom[25739] = 8'h06 ;
            rom[25740] = 8'hf5 ;
            rom[25741] = 8'h01 ;
            rom[25742] = 8'hfb ;
            rom[25743] = 8'he6 ;
            rom[25744] = 8'h07 ;
            rom[25745] = 8'h16 ;
            rom[25746] = 8'he6 ;
            rom[25747] = 8'hfb ;
            rom[25748] = 8'hd9 ;
            rom[25749] = 8'h19 ;
            rom[25750] = 8'hfc ;
            rom[25751] = 8'h08 ;
            rom[25752] = 8'hcc ;
            rom[25753] = 8'he3 ;
            rom[25754] = 8'h0f ;
            rom[25755] = 8'hc9 ;
            rom[25756] = 8'hf4 ;
            rom[25757] = 8'hd5 ;
            rom[25758] = 8'hbd ;
            rom[25759] = 8'h17 ;
            rom[25760] = 8'h16 ;
            rom[25761] = 8'h23 ;
            rom[25762] = 8'hf9 ;
            rom[25763] = 8'hf7 ;
            rom[25764] = 8'hed ;
            rom[25765] = 8'h0b ;
            rom[25766] = 8'h0b ;
            rom[25767] = 8'hc6 ;
            rom[25768] = 8'h05 ;
            rom[25769] = 8'h19 ;
            rom[25770] = 8'heb ;
            rom[25771] = 8'hf3 ;
            rom[25772] = 8'hd3 ;
            rom[25773] = 8'h15 ;
            rom[25774] = 8'h05 ;
            rom[25775] = 8'he0 ;
            rom[25776] = 8'he8 ;
            rom[25777] = 8'hde ;
            rom[25778] = 8'h1a ;
            rom[25779] = 8'h08 ;
            rom[25780] = 8'h0c ;
            rom[25781] = 8'hbc ;
            rom[25782] = 8'hfa ;
            rom[25783] = 8'h15 ;
            rom[25784] = 8'he2 ;
            rom[25785] = 8'hde ;
            rom[25786] = 8'hdb ;
            rom[25787] = 8'hf5 ;
            rom[25788] = 8'h0d ;
            rom[25789] = 8'h03 ;
            rom[25790] = 8'h08 ;
            rom[25791] = 8'hfb ;
            rom[25792] = 8'h19 ;
            rom[25793] = 8'he1 ;
            rom[25794] = 8'hec ;
            rom[25795] = 8'he1 ;
            rom[25796] = 8'hf0 ;
            rom[25797] = 8'h2c ;
            rom[25798] = 8'hed ;
            rom[25799] = 8'h17 ;
            rom[25800] = 8'h02 ;
            rom[25801] = 8'hfd ;
            rom[25802] = 8'h0d ;
            rom[25803] = 8'h1e ;
            rom[25804] = 8'he8 ;
            rom[25805] = 8'h00 ;
            rom[25806] = 8'h17 ;
            rom[25807] = 8'h12 ;
            rom[25808] = 8'hc0 ;
            rom[25809] = 8'h02 ;
            rom[25810] = 8'hfc ;
            rom[25811] = 8'h18 ;
            rom[25812] = 8'h0d ;
            rom[25813] = 8'hd0 ;
            rom[25814] = 8'hec ;
            rom[25815] = 8'hfa ;
            rom[25816] = 8'he8 ;
            rom[25817] = 8'hec ;
            rom[25818] = 8'h10 ;
            rom[25819] = 8'hfb ;
            rom[25820] = 8'hfd ;
            rom[25821] = 8'h08 ;
            rom[25822] = 8'hce ;
            rom[25823] = 8'h15 ;
            rom[25824] = 8'hec ;
            rom[25825] = 8'hfa ;
            rom[25826] = 8'h14 ;
            rom[25827] = 8'h03 ;
            rom[25828] = 8'hf5 ;
            rom[25829] = 8'hdc ;
            rom[25830] = 8'hf1 ;
            rom[25831] = 8'hf3 ;
            rom[25832] = 8'h11 ;
            rom[25833] = 8'hff ;
            rom[25834] = 8'hcf ;
            rom[25835] = 8'h03 ;
            rom[25836] = 8'hfa ;
            rom[25837] = 8'h16 ;
            rom[25838] = 8'h1d ;
            rom[25839] = 8'h08 ;
            rom[25840] = 8'hfb ;
            rom[25841] = 8'h1e ;
            rom[25842] = 8'h03 ;
            rom[25843] = 8'h0b ;
            rom[25844] = 8'h13 ;
            rom[25845] = 8'hf5 ;
            rom[25846] = 8'h0a ;
            rom[25847] = 8'h10 ;
            rom[25848] = 8'h09 ;
            rom[25849] = 8'hcc ;
            rom[25850] = 8'h0c ;
            rom[25851] = 8'h17 ;
            rom[25852] = 8'hf0 ;
            rom[25853] = 8'h21 ;
            rom[25854] = 8'he4 ;
            rom[25855] = 8'h12 ;
            rom[25856] = 8'h09 ;
            rom[25857] = 8'he5 ;
            rom[25858] = 8'hd5 ;
            rom[25859] = 8'hfa ;
            rom[25860] = 8'hf2 ;
            rom[25861] = 8'heb ;
            rom[25862] = 8'h1e ;
            rom[25863] = 8'hf9 ;
            rom[25864] = 8'hd6 ;
            rom[25865] = 8'h0e ;
            rom[25866] = 8'h05 ;
            rom[25867] = 8'h08 ;
            rom[25868] = 8'heb ;
            rom[25869] = 8'h0a ;
            rom[25870] = 8'h1f ;
            rom[25871] = 8'hf7 ;
            rom[25872] = 8'he2 ;
            rom[25873] = 8'h05 ;
            rom[25874] = 8'h05 ;
            rom[25875] = 8'hf7 ;
            rom[25876] = 8'h02 ;
            rom[25877] = 8'hdc ;
            rom[25878] = 8'hf5 ;
            rom[25879] = 8'hd9 ;
            rom[25880] = 8'he0 ;
            rom[25881] = 8'h17 ;
            rom[25882] = 8'h10 ;
            rom[25883] = 8'h19 ;
            rom[25884] = 8'h1b ;
            rom[25885] = 8'h13 ;
            rom[25886] = 8'hf7 ;
            rom[25887] = 8'h0f ;
            rom[25888] = 8'hfe ;
            rom[25889] = 8'he8 ;
            rom[25890] = 8'he9 ;
            rom[25891] = 8'h12 ;
            rom[25892] = 8'h08 ;
            rom[25893] = 8'hdf ;
            rom[25894] = 8'hdd ;
            rom[25895] = 8'heb ;
            rom[25896] = 8'h10 ;
            rom[25897] = 8'h0e ;
            rom[25898] = 8'h09 ;
            rom[25899] = 8'hd0 ;
            rom[25900] = 8'h06 ;
            rom[25901] = 8'he7 ;
            rom[25902] = 8'hcd ;
            rom[25903] = 8'hfe ;
            rom[25904] = 8'hed ;
            rom[25905] = 8'hff ;
            rom[25906] = 8'h31 ;
            rom[25907] = 8'hf1 ;
            rom[25908] = 8'hc4 ;
            rom[25909] = 8'he7 ;
            rom[25910] = 8'h11 ;
            rom[25911] = 8'h08 ;
            rom[25912] = 8'h0e ;
            rom[25913] = 8'h29 ;
            rom[25914] = 8'he4 ;
            rom[25915] = 8'h0f ;
            rom[25916] = 8'h0c ;
            rom[25917] = 8'hfb ;
            rom[25918] = 8'h01 ;
            rom[25919] = 8'hff ;
            rom[25920] = 8'h11 ;
            rom[25921] = 8'hde ;
            rom[25922] = 8'h1b ;
            rom[25923] = 8'hc6 ;
            rom[25924] = 8'hda ;
            rom[25925] = 8'h08 ;
            rom[25926] = 8'hca ;
            rom[25927] = 8'he5 ;
            rom[25928] = 8'h1d ;
            rom[25929] = 8'h01 ;
            rom[25930] = 8'h06 ;
            rom[25931] = 8'h14 ;
            rom[25932] = 8'he0 ;
            rom[25933] = 8'h2f ;
            rom[25934] = 8'h14 ;
            rom[25935] = 8'h20 ;
            rom[25936] = 8'h07 ;
            rom[25937] = 8'h01 ;
            rom[25938] = 8'hc7 ;
            rom[25939] = 8'hed ;
            rom[25940] = 8'h1d ;
            rom[25941] = 8'hc1 ;
            rom[25942] = 8'hdc ;
            rom[25943] = 8'hfc ;
            rom[25944] = 8'hd5 ;
            rom[25945] = 8'hcf ;
            rom[25946] = 8'hcc ;
            rom[25947] = 8'hf1 ;
            rom[25948] = 8'hf1 ;
            rom[25949] = 8'hf1 ;
            rom[25950] = 8'he4 ;
            rom[25951] = 8'h01 ;
            rom[25952] = 8'h1b ;
            rom[25953] = 8'h06 ;
            rom[25954] = 8'h19 ;
            rom[25955] = 8'hfc ;
            rom[25956] = 8'h0a ;
            rom[25957] = 8'hed ;
            rom[25958] = 8'h10 ;
            rom[25959] = 8'hfc ;
            rom[25960] = 8'hef ;
            rom[25961] = 8'h04 ;
            rom[25962] = 8'he2 ;
            rom[25963] = 8'h11 ;
            rom[25964] = 8'he6 ;
            rom[25965] = 8'h0a ;
            rom[25966] = 8'h00 ;
            rom[25967] = 8'hde ;
            rom[25968] = 8'hf4 ;
            rom[25969] = 8'h07 ;
            rom[25970] = 8'hec ;
            rom[25971] = 8'hf5 ;
            rom[25972] = 8'h11 ;
            rom[25973] = 8'hfa ;
            rom[25974] = 8'hd8 ;
            rom[25975] = 8'h25 ;
            rom[25976] = 8'h15 ;
            rom[25977] = 8'hff ;
            rom[25978] = 8'he9 ;
            rom[25979] = 8'hfc ;
            rom[25980] = 8'h06 ;
            rom[25981] = 8'h07 ;
            rom[25982] = 8'hfe ;
            rom[25983] = 8'hdc ;
            rom[25984] = 8'h23 ;
            rom[25985] = 8'h03 ;
            rom[25986] = 8'hf8 ;
            rom[25987] = 8'hed ;
            rom[25988] = 8'h18 ;
            rom[25989] = 8'hfa ;
            rom[25990] = 8'hec ;
            rom[25991] = 8'h18 ;
            rom[25992] = 8'hf0 ;
            rom[25993] = 8'he7 ;
            rom[25994] = 8'h06 ;
            rom[25995] = 8'hb6 ;
            rom[25996] = 8'hf6 ;
            rom[25997] = 8'he6 ;
            rom[25998] = 8'h10 ;
            rom[25999] = 8'hf1 ;
            rom[26000] = 8'h1d ;
            rom[26001] = 8'h04 ;
            rom[26002] = 8'h0e ;
            rom[26003] = 8'h06 ;
            rom[26004] = 8'hdb ;
            rom[26005] = 8'hbf ;
            rom[26006] = 8'hfa ;
            rom[26007] = 8'he8 ;
            rom[26008] = 8'hc4 ;
            rom[26009] = 8'hea ;
            rom[26010] = 8'hee ;
            rom[26011] = 8'hd6 ;
            rom[26012] = 8'h1a ;
            rom[26013] = 8'h00 ;
            rom[26014] = 8'h07 ;
            rom[26015] = 8'he9 ;
            rom[26016] = 8'h0f ;
            rom[26017] = 8'h29 ;
            rom[26018] = 8'h04 ;
            rom[26019] = 8'h22 ;
            rom[26020] = 8'hfc ;
            rom[26021] = 8'hef ;
            rom[26022] = 8'hca ;
            rom[26023] = 8'hfc ;
            rom[26024] = 8'hdb ;
            rom[26025] = 8'h08 ;
            rom[26026] = 8'hf6 ;
            rom[26027] = 8'h15 ;
            rom[26028] = 8'hf5 ;
            rom[26029] = 8'hbf ;
            rom[26030] = 8'hee ;
            rom[26031] = 8'h0b ;
            rom[26032] = 8'h1e ;
            rom[26033] = 8'hde ;
            rom[26034] = 8'hdc ;
            rom[26035] = 8'h11 ;
            rom[26036] = 8'hc8 ;
            rom[26037] = 8'h06 ;
            rom[26038] = 8'h1e ;
            rom[26039] = 8'hf7 ;
            rom[26040] = 8'hec ;
            rom[26041] = 8'h03 ;
            rom[26042] = 8'h27 ;
            rom[26043] = 8'hfe ;
            rom[26044] = 8'hf5 ;
            rom[26045] = 8'hf5 ;
            rom[26046] = 8'h25 ;
            rom[26047] = 8'he8 ;
            rom[26048] = 8'hef ;
            rom[26049] = 8'h08 ;
            rom[26050] = 8'he7 ;
            rom[26051] = 8'h0e ;
            rom[26052] = 8'hd1 ;
            rom[26053] = 8'h17 ;
            rom[26054] = 8'hfd ;
            rom[26055] = 8'h15 ;
            rom[26056] = 8'hfa ;
            rom[26057] = 8'h04 ;
            rom[26058] = 8'h00 ;
            rom[26059] = 8'hf3 ;
            rom[26060] = 8'hd0 ;
            rom[26061] = 8'he8 ;
            rom[26062] = 8'hfe ;
            rom[26063] = 8'hce ;
            rom[26064] = 8'h01 ;
            rom[26065] = 8'hc5 ;
            rom[26066] = 8'h08 ;
            rom[26067] = 8'hd3 ;
            rom[26068] = 8'h1a ;
            rom[26069] = 8'h04 ;
            rom[26070] = 8'hd0 ;
            rom[26071] = 8'hf6 ;
            rom[26072] = 8'hfc ;
            rom[26073] = 8'hd7 ;
            rom[26074] = 8'h0a ;
            rom[26075] = 8'h00 ;
            rom[26076] = 8'hfc ;
            rom[26077] = 8'hdf ;
            rom[26078] = 8'hf1 ;
            rom[26079] = 8'hfe ;
            rom[26080] = 8'hf6 ;
            rom[26081] = 8'hff ;
            rom[26082] = 8'hf9 ;
            rom[26083] = 8'h14 ;
            rom[26084] = 8'h0c ;
            rom[26085] = 8'h07 ;
            rom[26086] = 8'hfd ;
            rom[26087] = 8'h04 ;
            rom[26088] = 8'hcb ;
            rom[26089] = 8'h15 ;
            rom[26090] = 8'hf2 ;
            rom[26091] = 8'hf1 ;
            rom[26092] = 8'h01 ;
            rom[26093] = 8'h04 ;
            rom[26094] = 8'hef ;
            rom[26095] = 8'hd2 ;
            rom[26096] = 8'he5 ;
            rom[26097] = 8'hd5 ;
            rom[26098] = 8'hf7 ;
            rom[26099] = 8'h02 ;
            rom[26100] = 8'he4 ;
            rom[26101] = 8'hf1 ;
            rom[26102] = 8'hed ;
            rom[26103] = 8'h0f ;
            rom[26104] = 8'hf0 ;
            rom[26105] = 8'hcb ;
            rom[26106] = 8'hd4 ;
            rom[26107] = 8'hfb ;
            rom[26108] = 8'h04 ;
            rom[26109] = 8'hf2 ;
            rom[26110] = 8'h1a ;
            rom[26111] = 8'h15 ;
            rom[26112] = 8'hfc ;
            rom[26113] = 8'hc2 ;
            rom[26114] = 8'hfa ;
            rom[26115] = 8'hf4 ;
            rom[26116] = 8'hb4 ;
            rom[26117] = 8'hfe ;
            rom[26118] = 8'hf2 ;
            rom[26119] = 8'hf1 ;
            rom[26120] = 8'h0b ;
            rom[26121] = 8'h02 ;
            rom[26122] = 8'h0b ;
            rom[26123] = 8'hf9 ;
            rom[26124] = 8'h12 ;
            rom[26125] = 8'heb ;
            rom[26126] = 8'h00 ;
            rom[26127] = 8'he9 ;
            rom[26128] = 8'hfe ;
            rom[26129] = 8'he7 ;
            rom[26130] = 8'h0c ;
            rom[26131] = 8'h29 ;
            rom[26132] = 8'h03 ;
            rom[26133] = 8'he2 ;
            rom[26134] = 8'he7 ;
            rom[26135] = 8'h1b ;
            rom[26136] = 8'hd0 ;
            rom[26137] = 8'hfd ;
            rom[26138] = 8'hee ;
            rom[26139] = 8'hf6 ;
            rom[26140] = 8'h17 ;
            rom[26141] = 8'hf3 ;
            rom[26142] = 8'hea ;
            rom[26143] = 8'h07 ;
            rom[26144] = 8'hf8 ;
            rom[26145] = 8'hf7 ;
            rom[26146] = 8'h07 ;
            rom[26147] = 8'hcb ;
            rom[26148] = 8'h15 ;
            rom[26149] = 8'hf5 ;
            rom[26150] = 8'hff ;
            rom[26151] = 8'he4 ;
            rom[26152] = 8'hf2 ;
            rom[26153] = 8'he9 ;
            rom[26154] = 8'he9 ;
            rom[26155] = 8'hfc ;
            rom[26156] = 8'h19 ;
            rom[26157] = 8'hee ;
            rom[26158] = 8'heb ;
            rom[26159] = 8'hed ;
            rom[26160] = 8'h0a ;
            rom[26161] = 8'he6 ;
            rom[26162] = 8'h14 ;
            rom[26163] = 8'h28 ;
            rom[26164] = 8'he1 ;
            rom[26165] = 8'hfe ;
            rom[26166] = 8'hf2 ;
            rom[26167] = 8'hea ;
            rom[26168] = 8'h0a ;
            rom[26169] = 8'h18 ;
            rom[26170] = 8'hfd ;
            rom[26171] = 8'h01 ;
            rom[26172] = 8'he6 ;
            rom[26173] = 8'hfe ;
            rom[26174] = 8'h0e ;
            rom[26175] = 8'hfa ;
            rom[26176] = 8'h0e ;
            rom[26177] = 8'hfb ;
            rom[26178] = 8'h06 ;
            rom[26179] = 8'hfe ;
            rom[26180] = 8'h0f ;
            rom[26181] = 8'h36 ;
            rom[26182] = 8'h18 ;
            rom[26183] = 8'hdb ;
            rom[26184] = 8'hde ;
            rom[26185] = 8'hfc ;
            rom[26186] = 8'heb ;
            rom[26187] = 8'h1b ;
            rom[26188] = 8'hd5 ;
            rom[26189] = 8'h0b ;
            rom[26190] = 8'h09 ;
            rom[26191] = 8'hf6 ;
            rom[26192] = 8'h0c ;
            rom[26193] = 8'hf7 ;
            rom[26194] = 8'h0d ;
            rom[26195] = 8'hd4 ;
            rom[26196] = 8'h14 ;
            rom[26197] = 8'he2 ;
            rom[26198] = 8'hef ;
            rom[26199] = 8'hf0 ;
            rom[26200] = 8'hfe ;
            rom[26201] = 8'he0 ;
            rom[26202] = 8'hd9 ;
            rom[26203] = 8'he2 ;
            rom[26204] = 8'hef ;
            rom[26205] = 8'hda ;
            rom[26206] = 8'h07 ;
            rom[26207] = 8'hc9 ;
            rom[26208] = 8'hec ;
            rom[26209] = 8'hff ;
            rom[26210] = 8'hd4 ;
            rom[26211] = 8'h0d ;
            rom[26212] = 8'he4 ;
            rom[26213] = 8'hf0 ;
            rom[26214] = 8'h01 ;
            rom[26215] = 8'h02 ;
            rom[26216] = 8'h0f ;
            rom[26217] = 8'hf9 ;
            rom[26218] = 8'h00 ;
            rom[26219] = 8'h19 ;
            rom[26220] = 8'hf4 ;
            rom[26221] = 8'he8 ;
            rom[26222] = 8'hec ;
            rom[26223] = 8'hd1 ;
            rom[26224] = 8'h07 ;
            rom[26225] = 8'h11 ;
            rom[26226] = 8'hf7 ;
            rom[26227] = 8'hd9 ;
            rom[26228] = 8'h1a ;
            rom[26229] = 8'he9 ;
            rom[26230] = 8'he8 ;
            rom[26231] = 8'h06 ;
            rom[26232] = 8'hf4 ;
            rom[26233] = 8'he8 ;
            rom[26234] = 8'hd7 ;
            rom[26235] = 8'hf3 ;
            rom[26236] = 8'h0b ;
            rom[26237] = 8'h2e ;
            rom[26238] = 8'hd5 ;
            rom[26239] = 8'h07 ;
            rom[26240] = 8'hcf ;
            rom[26241] = 8'hd8 ;
            rom[26242] = 8'hf9 ;
            rom[26243] = 8'h0e ;
            rom[26244] = 8'h3d ;
            rom[26245] = 8'h02 ;
            rom[26246] = 8'h10 ;
            rom[26247] = 8'h19 ;
            rom[26248] = 8'he6 ;
            rom[26249] = 8'h0d ;
            rom[26250] = 8'h16 ;
            rom[26251] = 8'hfc ;
            rom[26252] = 8'h04 ;
            rom[26253] = 8'hea ;
            rom[26254] = 8'h09 ;
            rom[26255] = 8'h09 ;
            rom[26256] = 8'h05 ;
            rom[26257] = 8'he8 ;
            rom[26258] = 8'h08 ;
            rom[26259] = 8'h0d ;
            rom[26260] = 8'hf2 ;
            rom[26261] = 8'h0a ;
            rom[26262] = 8'h10 ;
            rom[26263] = 8'h09 ;
            rom[26264] = 8'he9 ;
            rom[26265] = 8'hcb ;
            rom[26266] = 8'h20 ;
            rom[26267] = 8'hfe ;
            rom[26268] = 8'hf9 ;
            rom[26269] = 8'hef ;
            rom[26270] = 8'h14 ;
            rom[26271] = 8'h0a ;
            rom[26272] = 8'h25 ;
            rom[26273] = 8'h07 ;
            rom[26274] = 8'hde ;
            rom[26275] = 8'h03 ;
            rom[26276] = 8'hf1 ;
            rom[26277] = 8'hf1 ;
            rom[26278] = 8'hf0 ;
            rom[26279] = 8'hfc ;
            rom[26280] = 8'hdf ;
            rom[26281] = 8'hea ;
            rom[26282] = 8'hf9 ;
            rom[26283] = 8'h11 ;
            rom[26284] = 8'h0b ;
            rom[26285] = 8'hd5 ;
            rom[26286] = 8'hf1 ;
            rom[26287] = 8'hf4 ;
            rom[26288] = 8'hf6 ;
            rom[26289] = 8'h11 ;
            rom[26290] = 8'h03 ;
            rom[26291] = 8'hd6 ;
            rom[26292] = 8'hcb ;
            rom[26293] = 8'hfe ;
            rom[26294] = 8'h39 ;
            rom[26295] = 8'hf3 ;
            rom[26296] = 8'hd0 ;
            rom[26297] = 8'hf7 ;
            rom[26298] = 8'h08 ;
            rom[26299] = 8'h1d ;
            rom[26300] = 8'hec ;
            rom[26301] = 8'h15 ;
            rom[26302] = 8'hfb ;
            rom[26303] = 8'h01 ;
            rom[26304] = 8'h06 ;
            rom[26305] = 8'hdf ;
            rom[26306] = 8'he7 ;
            rom[26307] = 8'hc4 ;
            rom[26308] = 8'he7 ;
            rom[26309] = 8'hdf ;
            rom[26310] = 8'hf1 ;
            rom[26311] = 8'h0f ;
            rom[26312] = 8'h01 ;
            rom[26313] = 8'h06 ;
            rom[26314] = 8'h1c ;
            rom[26315] = 8'h28 ;
            rom[26316] = 8'hff ;
            rom[26317] = 8'hfb ;
            rom[26318] = 8'hfe ;
            rom[26319] = 8'h01 ;
            rom[26320] = 8'hd8 ;
            rom[26321] = 8'h11 ;
            rom[26322] = 8'hf9 ;
            rom[26323] = 8'h08 ;
            rom[26324] = 8'h0a ;
            rom[26325] = 8'hed ;
            rom[26326] = 8'h12 ;
            rom[26327] = 8'hd2 ;
            rom[26328] = 8'he8 ;
            rom[26329] = 8'h1f ;
            rom[26330] = 8'h08 ;
            rom[26331] = 8'hfb ;
            rom[26332] = 8'h18 ;
            rom[26333] = 8'h09 ;
            rom[26334] = 8'h23 ;
            rom[26335] = 8'hf4 ;
            rom[26336] = 8'h10 ;
            rom[26337] = 8'h1a ;
            rom[26338] = 8'h0b ;
            rom[26339] = 8'hf6 ;
            rom[26340] = 8'hfa ;
            rom[26341] = 8'hd3 ;
            rom[26342] = 8'h04 ;
            rom[26343] = 8'h0a ;
            rom[26344] = 8'h08 ;
            rom[26345] = 8'hfa ;
            rom[26346] = 8'hbf ;
            rom[26347] = 8'hfc ;
            rom[26348] = 8'hf5 ;
            rom[26349] = 8'h18 ;
            rom[26350] = 8'h00 ;
            rom[26351] = 8'h0d ;
            rom[26352] = 8'h09 ;
            rom[26353] = 8'hfa ;
            rom[26354] = 8'hf1 ;
            rom[26355] = 8'hd2 ;
            rom[26356] = 8'h08 ;
            rom[26357] = 8'he9 ;
            rom[26358] = 8'he4 ;
            rom[26359] = 8'h00 ;
            rom[26360] = 8'h0e ;
            rom[26361] = 8'h17 ;
            rom[26362] = 8'hfc ;
            rom[26363] = 8'h05 ;
            rom[26364] = 8'hfb ;
            rom[26365] = 8'hfa ;
            rom[26366] = 8'hf6 ;
            rom[26367] = 8'h00 ;
            rom[26368] = 8'hfc ;
            rom[26369] = 8'h04 ;
            rom[26370] = 8'h22 ;
            rom[26371] = 8'h2d ;
            rom[26372] = 8'h04 ;
            rom[26373] = 8'h00 ;
            rom[26374] = 8'hec ;
            rom[26375] = 8'he8 ;
            rom[26376] = 8'he4 ;
            rom[26377] = 8'h02 ;
            rom[26378] = 8'h00 ;
            rom[26379] = 8'hdc ;
            rom[26380] = 8'h09 ;
            rom[26381] = 8'hfe ;
            rom[26382] = 8'h20 ;
            rom[26383] = 8'h19 ;
            rom[26384] = 8'h11 ;
            rom[26385] = 8'h0b ;
            rom[26386] = 8'h13 ;
            rom[26387] = 8'h13 ;
            rom[26388] = 8'he8 ;
            rom[26389] = 8'hca ;
            rom[26390] = 8'hfd ;
            rom[26391] = 8'h13 ;
            rom[26392] = 8'hf5 ;
            rom[26393] = 8'he0 ;
            rom[26394] = 8'h00 ;
            rom[26395] = 8'he6 ;
            rom[26396] = 8'hda ;
            rom[26397] = 8'hea ;
            rom[26398] = 8'hff ;
            rom[26399] = 8'hda ;
            rom[26400] = 8'h0a ;
            rom[26401] = 8'h34 ;
            rom[26402] = 8'he6 ;
            rom[26403] = 8'hf5 ;
            rom[26404] = 8'h06 ;
            rom[26405] = 8'h0a ;
            rom[26406] = 8'he4 ;
            rom[26407] = 8'hfe ;
            rom[26408] = 8'hf3 ;
            rom[26409] = 8'hc1 ;
            rom[26410] = 8'h0a ;
            rom[26411] = 8'h0a ;
            rom[26412] = 8'hdc ;
            rom[26413] = 8'hf1 ;
            rom[26414] = 8'h18 ;
            rom[26415] = 8'hf4 ;
            rom[26416] = 8'hfd ;
            rom[26417] = 8'h02 ;
            rom[26418] = 8'hd9 ;
            rom[26419] = 8'hf4 ;
            rom[26420] = 8'h10 ;
            rom[26421] = 8'h0e ;
            rom[26422] = 8'hff ;
            rom[26423] = 8'hda ;
            rom[26424] = 8'h16 ;
            rom[26425] = 8'h16 ;
            rom[26426] = 8'h08 ;
            rom[26427] = 8'hdb ;
            rom[26428] = 8'hf9 ;
            rom[26429] = 8'hf6 ;
            rom[26430] = 8'hfc ;
            rom[26431] = 8'h0c ;
            rom[26432] = 8'hdb ;
            rom[26433] = 8'hfb ;
            rom[26434] = 8'h10 ;
            rom[26435] = 8'h08 ;
            rom[26436] = 8'hcc ;
            rom[26437] = 8'h15 ;
            rom[26438] = 8'hd7 ;
            rom[26439] = 8'hf1 ;
            rom[26440] = 8'he9 ;
            rom[26441] = 8'hfa ;
            rom[26442] = 8'h1f ;
            rom[26443] = 8'hea ;
            rom[26444] = 8'h0a ;
            rom[26445] = 8'h16 ;
            rom[26446] = 8'hed ;
            rom[26447] = 8'h09 ;
            rom[26448] = 8'h0e ;
            rom[26449] = 8'hf8 ;
            rom[26450] = 8'hfc ;
            rom[26451] = 8'h0d ;
            rom[26452] = 8'h0e ;
            rom[26453] = 8'hde ;
            rom[26454] = 8'hff ;
            rom[26455] = 8'h08 ;
            rom[26456] = 8'h0e ;
            rom[26457] = 8'h04 ;
            rom[26458] = 8'h1b ;
            rom[26459] = 8'h13 ;
            rom[26460] = 8'h11 ;
            rom[26461] = 8'hf8 ;
            rom[26462] = 8'h01 ;
            rom[26463] = 8'h16 ;
            rom[26464] = 8'h19 ;
            rom[26465] = 8'he2 ;
            rom[26466] = 8'hff ;
            rom[26467] = 8'hfd ;
            rom[26468] = 8'he4 ;
            rom[26469] = 8'hf5 ;
            rom[26470] = 8'h17 ;
            rom[26471] = 8'h03 ;
            rom[26472] = 8'he2 ;
            rom[26473] = 8'hf2 ;
            rom[26474] = 8'h00 ;
            rom[26475] = 8'hf1 ;
            rom[26476] = 8'h13 ;
            rom[26477] = 8'h04 ;
            rom[26478] = 8'h12 ;
            rom[26479] = 8'h00 ;
            rom[26480] = 8'h2f ;
            rom[26481] = 8'hdb ;
            rom[26482] = 8'h03 ;
            rom[26483] = 8'heb ;
            rom[26484] = 8'hef ;
            rom[26485] = 8'h07 ;
            rom[26486] = 8'hc4 ;
            rom[26487] = 8'hf8 ;
            rom[26488] = 8'he7 ;
            rom[26489] = 8'h07 ;
            rom[26490] = 8'h1a ;
            rom[26491] = 8'hbe ;
            rom[26492] = 8'hec ;
            rom[26493] = 8'h01 ;
            rom[26494] = 8'he0 ;
            rom[26495] = 8'hea ;
            rom[26496] = 8'hfc ;
            rom[26497] = 8'hf3 ;
            rom[26498] = 8'h0d ;
            rom[26499] = 8'h1a ;
            rom[26500] = 8'h0d ;
            rom[26501] = 8'h1b ;
            rom[26502] = 8'h32 ;
            rom[26503] = 8'h11 ;
            rom[26504] = 8'h27 ;
            rom[26505] = 8'h13 ;
            rom[26506] = 8'hdb ;
            rom[26507] = 8'hfc ;
            rom[26508] = 8'h06 ;
            rom[26509] = 8'hfb ;
            rom[26510] = 8'hf3 ;
            rom[26511] = 8'h2a ;
            rom[26512] = 8'hf0 ;
            rom[26513] = 8'hd4 ;
            rom[26514] = 8'h09 ;
            rom[26515] = 8'h19 ;
            rom[26516] = 8'h23 ;
            rom[26517] = 8'hf5 ;
            rom[26518] = 8'h03 ;
            rom[26519] = 8'h12 ;
            rom[26520] = 8'h0c ;
            rom[26521] = 8'h0b ;
            rom[26522] = 8'h0e ;
            rom[26523] = 8'hdd ;
            rom[26524] = 8'hf5 ;
            rom[26525] = 8'hf0 ;
            rom[26526] = 8'h2c ;
            rom[26527] = 8'h0c ;
            rom[26528] = 8'h1b ;
            rom[26529] = 8'h06 ;
            rom[26530] = 8'hf2 ;
            rom[26531] = 8'h04 ;
            rom[26532] = 8'h17 ;
            rom[26533] = 8'h25 ;
            rom[26534] = 8'hff ;
            rom[26535] = 8'hf8 ;
            rom[26536] = 8'hdc ;
            rom[26537] = 8'he1 ;
            rom[26538] = 8'hf9 ;
            rom[26539] = 8'hee ;
            rom[26540] = 8'h05 ;
            rom[26541] = 8'h0e ;
            rom[26542] = 8'he5 ;
            rom[26543] = 8'h0b ;
            rom[26544] = 8'hf6 ;
            rom[26545] = 8'h1d ;
            rom[26546] = 8'hfc ;
            rom[26547] = 8'hfd ;
            rom[26548] = 8'hf7 ;
            rom[26549] = 8'hf4 ;
            rom[26550] = 8'he8 ;
            rom[26551] = 8'hd6 ;
            rom[26552] = 8'h0d ;
            rom[26553] = 8'h0b ;
            rom[26554] = 8'h19 ;
            rom[26555] = 8'hfd ;
            rom[26556] = 8'hea ;
            rom[26557] = 8'hfb ;
            rom[26558] = 8'hd9 ;
            rom[26559] = 8'he9 ;
            rom[26560] = 8'h06 ;
            rom[26561] = 8'h0a ;
            rom[26562] = 8'h25 ;
            rom[26563] = 8'he3 ;
            rom[26564] = 8'hf1 ;
            rom[26565] = 8'hdc ;
            rom[26566] = 8'hf2 ;
            rom[26567] = 8'hc0 ;
            rom[26568] = 8'h0d ;
            rom[26569] = 8'hd3 ;
            rom[26570] = 8'h22 ;
            rom[26571] = 8'hea ;
            rom[26572] = 8'hfb ;
            rom[26573] = 8'hee ;
            rom[26574] = 8'hf7 ;
            rom[26575] = 8'h04 ;
            rom[26576] = 8'h14 ;
            rom[26577] = 8'h05 ;
            rom[26578] = 8'hed ;
            rom[26579] = 8'h1f ;
            rom[26580] = 8'hd6 ;
            rom[26581] = 8'hd1 ;
            rom[26582] = 8'h26 ;
            rom[26583] = 8'hd1 ;
            rom[26584] = 8'hdb ;
            rom[26585] = 8'hec ;
            rom[26586] = 8'h10 ;
            rom[26587] = 8'h26 ;
            rom[26588] = 8'hf8 ;
            rom[26589] = 8'hfa ;
            rom[26590] = 8'hee ;
            rom[26591] = 8'h06 ;
            rom[26592] = 8'h13 ;
            rom[26593] = 8'hfe ;
            rom[26594] = 8'hdf ;
            rom[26595] = 8'h10 ;
            rom[26596] = 8'h1f ;
            rom[26597] = 8'he3 ;
            rom[26598] = 8'h02 ;
            rom[26599] = 8'hdd ;
            rom[26600] = 8'hf3 ;
            rom[26601] = 8'he5 ;
            rom[26602] = 8'hfe ;
            rom[26603] = 8'h26 ;
            rom[26604] = 8'he6 ;
            rom[26605] = 8'he6 ;
            rom[26606] = 8'h01 ;
            rom[26607] = 8'heb ;
            rom[26608] = 8'h10 ;
            rom[26609] = 8'he3 ;
            rom[26610] = 8'hfd ;
            rom[26611] = 8'hfd ;
            rom[26612] = 8'he5 ;
            rom[26613] = 8'hd3 ;
            rom[26614] = 8'hfa ;
            rom[26615] = 8'hd9 ;
            rom[26616] = 8'hd2 ;
            rom[26617] = 8'h03 ;
            rom[26618] = 8'h0a ;
            rom[26619] = 8'h0b ;
            rom[26620] = 8'hd9 ;
            rom[26621] = 8'hd0 ;
            rom[26622] = 8'hef ;
            rom[26623] = 8'h0a ;
            rom[26624] = 8'hf8 ;
            rom[26625] = 8'hfc ;
            rom[26626] = 8'h09 ;
            rom[26627] = 8'h14 ;
            rom[26628] = 8'h15 ;
            rom[26629] = 8'h02 ;
            rom[26630] = 8'h0f ;
            rom[26631] = 8'h0b ;
            rom[26632] = 8'hf5 ;
            rom[26633] = 8'h2b ;
            rom[26634] = 8'hf4 ;
            rom[26635] = 8'h14 ;
            rom[26636] = 8'hef ;
            rom[26637] = 8'h10 ;
            rom[26638] = 8'hcd ;
            rom[26639] = 8'hfe ;
            rom[26640] = 8'h03 ;
            rom[26641] = 8'h0c ;
            rom[26642] = 8'hf4 ;
            rom[26643] = 8'h04 ;
            rom[26644] = 8'h11 ;
            rom[26645] = 8'h0a ;
            rom[26646] = 8'hff ;
            rom[26647] = 8'hf5 ;
            rom[26648] = 8'h11 ;
            rom[26649] = 8'h33 ;
            rom[26650] = 8'h15 ;
            rom[26651] = 8'h28 ;
            rom[26652] = 8'h10 ;
            rom[26653] = 8'he0 ;
            rom[26654] = 8'h2e ;
            rom[26655] = 8'h1f ;
            rom[26656] = 8'h1c ;
            rom[26657] = 8'h03 ;
            rom[26658] = 8'hd3 ;
            rom[26659] = 8'h06 ;
            rom[26660] = 8'h02 ;
            rom[26661] = 8'hec ;
            rom[26662] = 8'h04 ;
            rom[26663] = 8'h1c ;
            rom[26664] = 8'h27 ;
            rom[26665] = 8'h06 ;
            rom[26666] = 8'hf1 ;
            rom[26667] = 8'h17 ;
            rom[26668] = 8'h04 ;
            rom[26669] = 8'hf2 ;
            rom[26670] = 8'h02 ;
            rom[26671] = 8'he8 ;
            rom[26672] = 8'hfb ;
            rom[26673] = 8'h0f ;
            rom[26674] = 8'h16 ;
            rom[26675] = 8'h08 ;
            rom[26676] = 8'hcd ;
            rom[26677] = 8'he5 ;
            rom[26678] = 8'h13 ;
            rom[26679] = 8'h02 ;
            rom[26680] = 8'hf2 ;
            rom[26681] = 8'h08 ;
            rom[26682] = 8'h14 ;
            rom[26683] = 8'h1e ;
            rom[26684] = 8'hef ;
            rom[26685] = 8'h25 ;
            rom[26686] = 8'hd7 ;
            rom[26687] = 8'h16 ;
            rom[26688] = 8'h0c ;
            rom[26689] = 8'he6 ;
            rom[26690] = 8'hfa ;
            rom[26691] = 8'hbd ;
            rom[26692] = 8'hee ;
            rom[26693] = 8'hc3 ;
            rom[26694] = 8'h0a ;
            rom[26695] = 8'hca ;
            rom[26696] = 8'hfb ;
            rom[26697] = 8'hfc ;
            rom[26698] = 8'h18 ;
            rom[26699] = 8'h14 ;
            rom[26700] = 8'h08 ;
            rom[26701] = 8'h1f ;
            rom[26702] = 8'h12 ;
            rom[26703] = 8'h25 ;
            rom[26704] = 8'h03 ;
            rom[26705] = 8'h00 ;
            rom[26706] = 8'hcb ;
            rom[26707] = 8'he8 ;
            rom[26708] = 8'h20 ;
            rom[26709] = 8'ha1 ;
            rom[26710] = 8'hfa ;
            rom[26711] = 8'hde ;
            rom[26712] = 8'h16 ;
            rom[26713] = 8'h19 ;
            rom[26714] = 8'hd9 ;
            rom[26715] = 8'h05 ;
            rom[26716] = 8'h06 ;
            rom[26717] = 8'h17 ;
            rom[26718] = 8'h08 ;
            rom[26719] = 8'hde ;
            rom[26720] = 8'h06 ;
            rom[26721] = 8'hff ;
            rom[26722] = 8'he3 ;
            rom[26723] = 8'hfb ;
            rom[26724] = 8'h21 ;
            rom[26725] = 8'hf7 ;
            rom[26726] = 8'hdf ;
            rom[26727] = 8'h20 ;
            rom[26728] = 8'hf1 ;
            rom[26729] = 8'h01 ;
            rom[26730] = 8'he4 ;
            rom[26731] = 8'hfb ;
            rom[26732] = 8'h89 ;
            rom[26733] = 8'hda ;
            rom[26734] = 8'hdc ;
            rom[26735] = 8'h13 ;
            rom[26736] = 8'h22 ;
            rom[26737] = 8'h1b ;
            rom[26738] = 8'h20 ;
            rom[26739] = 8'hd4 ;
            rom[26740] = 8'h13 ;
            rom[26741] = 8'h08 ;
            rom[26742] = 8'hfb ;
            rom[26743] = 8'hfc ;
            rom[26744] = 8'h04 ;
            rom[26745] = 8'h10 ;
            rom[26746] = 8'h00 ;
            rom[26747] = 8'h37 ;
            rom[26748] = 8'hdc ;
            rom[26749] = 8'he4 ;
            rom[26750] = 8'hd9 ;
            rom[26751] = 8'h0a ;
            rom[26752] = 8'h21 ;
            rom[26753] = 8'h02 ;
            rom[26754] = 8'h12 ;
            rom[26755] = 8'hf5 ;
            rom[26756] = 8'hfb ;
            rom[26757] = 8'h0a ;
            rom[26758] = 8'h1e ;
            rom[26759] = 8'h0e ;
            rom[26760] = 8'h08 ;
            rom[26761] = 8'hde ;
            rom[26762] = 8'hee ;
            rom[26763] = 8'he6 ;
            rom[26764] = 8'h0b ;
            rom[26765] = 8'he0 ;
            rom[26766] = 8'hfd ;
            rom[26767] = 8'hc8 ;
            rom[26768] = 8'hf6 ;
            rom[26769] = 8'h0e ;
            rom[26770] = 8'h21 ;
            rom[26771] = 8'h09 ;
            rom[26772] = 8'hed ;
            rom[26773] = 8'hd6 ;
            rom[26774] = 8'h00 ;
            rom[26775] = 8'hd5 ;
            rom[26776] = 8'hd2 ;
            rom[26777] = 8'h12 ;
            rom[26778] = 8'hce ;
            rom[26779] = 8'hf2 ;
            rom[26780] = 8'h03 ;
            rom[26781] = 8'hff ;
            rom[26782] = 8'hf2 ;
            rom[26783] = 8'h09 ;
            rom[26784] = 8'he7 ;
            rom[26785] = 8'h05 ;
            rom[26786] = 8'h03 ;
            rom[26787] = 8'hef ;
            rom[26788] = 8'h0f ;
            rom[26789] = 8'h0c ;
            rom[26790] = 8'h2c ;
            rom[26791] = 8'hec ;
            rom[26792] = 8'hee ;
            rom[26793] = 8'hdf ;
            rom[26794] = 8'h08 ;
            rom[26795] = 8'he4 ;
            rom[26796] = 8'h00 ;
            rom[26797] = 8'h0c ;
            rom[26798] = 8'hee ;
            rom[26799] = 8'h26 ;
            rom[26800] = 8'he3 ;
            rom[26801] = 8'h05 ;
            rom[26802] = 8'h13 ;
            rom[26803] = 8'h25 ;
            rom[26804] = 8'hd2 ;
            rom[26805] = 8'hf1 ;
            rom[26806] = 8'hf2 ;
            rom[26807] = 8'h21 ;
            rom[26808] = 8'hcb ;
            rom[26809] = 8'h1b ;
            rom[26810] = 8'h25 ;
            rom[26811] = 8'hea ;
            rom[26812] = 8'hf9 ;
            rom[26813] = 8'h02 ;
            rom[26814] = 8'hf1 ;
            rom[26815] = 8'he8 ;
            rom[26816] = 8'he8 ;
            rom[26817] = 8'h24 ;
            rom[26818] = 8'hf2 ;
            rom[26819] = 8'h0a ;
            rom[26820] = 8'h0e ;
            rom[26821] = 8'h02 ;
            rom[26822] = 8'h00 ;
            rom[26823] = 8'h1c ;
            rom[26824] = 8'hd2 ;
            rom[26825] = 8'h12 ;
            rom[26826] = 8'hff ;
            rom[26827] = 8'hff ;
            rom[26828] = 8'h07 ;
            rom[26829] = 8'h03 ;
            rom[26830] = 8'hed ;
            rom[26831] = 8'hfd ;
            rom[26832] = 8'he4 ;
            rom[26833] = 8'h00 ;
            rom[26834] = 8'h2b ;
            rom[26835] = 8'hd1 ;
            rom[26836] = 8'hfa ;
            rom[26837] = 8'hfc ;
            rom[26838] = 8'h01 ;
            rom[26839] = 8'h23 ;
            rom[26840] = 8'h0d ;
            rom[26841] = 8'h25 ;
            rom[26842] = 8'h2c ;
            rom[26843] = 8'h08 ;
            rom[26844] = 8'hf2 ;
            rom[26845] = 8'hc8 ;
            rom[26846] = 8'hf6 ;
            rom[26847] = 8'hee ;
            rom[26848] = 8'hfc ;
            rom[26849] = 8'h2f ;
            rom[26850] = 8'hf6 ;
            rom[26851] = 8'h08 ;
            rom[26852] = 8'he5 ;
            rom[26853] = 8'he8 ;
            rom[26854] = 8'hff ;
            rom[26855] = 8'h0b ;
            rom[26856] = 8'h05 ;
            rom[26857] = 8'hf6 ;
            rom[26858] = 8'h1a ;
            rom[26859] = 8'he8 ;
            rom[26860] = 8'h07 ;
            rom[26861] = 8'h0f ;
            rom[26862] = 8'h00 ;
            rom[26863] = 8'hd0 ;
            rom[26864] = 8'hba ;
            rom[26865] = 8'h07 ;
            rom[26866] = 8'h07 ;
            rom[26867] = 8'h13 ;
            rom[26868] = 8'he3 ;
            rom[26869] = 8'hf9 ;
            rom[26870] = 8'hea ;
            rom[26871] = 8'h0d ;
            rom[26872] = 8'h13 ;
            rom[26873] = 8'he7 ;
            rom[26874] = 8'h07 ;
            rom[26875] = 8'h0a ;
            rom[26876] = 8'hd7 ;
            rom[26877] = 8'hf5 ;
            rom[26878] = 8'hf5 ;
            rom[26879] = 8'hdc ;
            rom[26880] = 8'h0d ;
            rom[26881] = 8'h0b ;
            rom[26882] = 8'he3 ;
            rom[26883] = 8'hdf ;
            rom[26884] = 8'hea ;
            rom[26885] = 8'h07 ;
            rom[26886] = 8'hf6 ;
            rom[26887] = 8'h0e ;
            rom[26888] = 8'h08 ;
            rom[26889] = 8'he0 ;
            rom[26890] = 8'hf3 ;
            rom[26891] = 8'h02 ;
            rom[26892] = 8'hec ;
            rom[26893] = 8'h0a ;
            rom[26894] = 8'h13 ;
            rom[26895] = 8'h17 ;
            rom[26896] = 8'hfc ;
            rom[26897] = 8'he1 ;
            rom[26898] = 8'hfb ;
            rom[26899] = 8'hf6 ;
            rom[26900] = 8'hec ;
            rom[26901] = 8'h08 ;
            rom[26902] = 8'h0e ;
            rom[26903] = 8'h06 ;
            rom[26904] = 8'he9 ;
            rom[26905] = 8'he2 ;
            rom[26906] = 8'hf9 ;
            rom[26907] = 8'h09 ;
            rom[26908] = 8'h1a ;
            rom[26909] = 8'hfb ;
            rom[26910] = 8'hf3 ;
            rom[26911] = 8'hbd ;
            rom[26912] = 8'hf3 ;
            rom[26913] = 8'h17 ;
            rom[26914] = 8'h09 ;
            rom[26915] = 8'h06 ;
            rom[26916] = 8'hff ;
            rom[26917] = 8'h23 ;
            rom[26918] = 8'he2 ;
            rom[26919] = 8'hd5 ;
            rom[26920] = 8'h13 ;
            rom[26921] = 8'hd4 ;
            rom[26922] = 8'h3a ;
            rom[26923] = 8'he1 ;
            rom[26924] = 8'hfd ;
            rom[26925] = 8'hfc ;
            rom[26926] = 8'h03 ;
            rom[26927] = 8'h06 ;
            rom[26928] = 8'he8 ;
            rom[26929] = 8'hf4 ;
            rom[26930] = 8'hf1 ;
            rom[26931] = 8'hc0 ;
            rom[26932] = 8'h09 ;
            rom[26933] = 8'hdb ;
            rom[26934] = 8'he4 ;
            rom[26935] = 8'h11 ;
            rom[26936] = 8'hfa ;
            rom[26937] = 8'h11 ;
            rom[26938] = 8'hf4 ;
            rom[26939] = 8'hd5 ;
            rom[26940] = 8'h08 ;
            rom[26941] = 8'h10 ;
            rom[26942] = 8'he4 ;
            rom[26943] = 8'hb8 ;
            rom[26944] = 8'h05 ;
            rom[26945] = 8'hec ;
            rom[26946] = 8'hf6 ;
            rom[26947] = 8'h21 ;
            rom[26948] = 8'hf1 ;
            rom[26949] = 8'hf5 ;
            rom[26950] = 8'he8 ;
            rom[26951] = 8'h00 ;
            rom[26952] = 8'h08 ;
            rom[26953] = 8'h0f ;
            rom[26954] = 8'hf1 ;
            rom[26955] = 8'h0b ;
            rom[26956] = 8'hf4 ;
            rom[26957] = 8'h04 ;
            rom[26958] = 8'h1f ;
            rom[26959] = 8'h3b ;
            rom[26960] = 8'hfc ;
            rom[26961] = 8'h1d ;
            rom[26962] = 8'h23 ;
            rom[26963] = 8'h18 ;
            rom[26964] = 8'h17 ;
            rom[26965] = 8'he3 ;
            rom[26966] = 8'h09 ;
            rom[26967] = 8'hf4 ;
            rom[26968] = 8'hf8 ;
            rom[26969] = 8'hed ;
            rom[26970] = 8'hed ;
            rom[26971] = 8'hfb ;
            rom[26972] = 8'he1 ;
            rom[26973] = 8'hfa ;
            rom[26974] = 8'he9 ;
            rom[26975] = 8'h21 ;
            rom[26976] = 8'h03 ;
            rom[26977] = 8'h17 ;
            rom[26978] = 8'h05 ;
            rom[26979] = 8'hd9 ;
            rom[26980] = 8'he9 ;
            rom[26981] = 8'hd7 ;
            rom[26982] = 8'he3 ;
            rom[26983] = 8'h17 ;
            rom[26984] = 8'h10 ;
            rom[26985] = 8'h04 ;
            rom[26986] = 8'hea ;
            rom[26987] = 8'h05 ;
            rom[26988] = 8'h05 ;
            rom[26989] = 8'h1d ;
            rom[26990] = 8'h08 ;
            rom[26991] = 8'hdb ;
            rom[26992] = 8'hf8 ;
            rom[26993] = 8'he3 ;
            rom[26994] = 8'h09 ;
            rom[26995] = 8'h1c ;
            rom[26996] = 8'hff ;
            rom[26997] = 8'h1d ;
            rom[26998] = 8'h06 ;
            rom[26999] = 8'h01 ;
            rom[27000] = 8'hff ;
            rom[27001] = 8'h12 ;
            rom[27002] = 8'hf7 ;
            rom[27003] = 8'he8 ;
            rom[27004] = 8'h05 ;
            rom[27005] = 8'he5 ;
            rom[27006] = 8'h05 ;
            rom[27007] = 8'h10 ;
            rom[27008] = 8'hf2 ;
            rom[27009] = 8'he5 ;
            rom[27010] = 8'he3 ;
            rom[27011] = 8'h25 ;
            rom[27012] = 8'hf5 ;
            rom[27013] = 8'hfc ;
            rom[27014] = 8'h22 ;
            rom[27015] = 8'h0b ;
            rom[27016] = 8'hf3 ;
            rom[27017] = 8'h46 ;
            rom[27018] = 8'hee ;
            rom[27019] = 8'hfa ;
            rom[27020] = 8'hfc ;
            rom[27021] = 8'hf9 ;
            rom[27022] = 8'he1 ;
            rom[27023] = 8'hf7 ;
            rom[27024] = 8'hed ;
            rom[27025] = 8'hf2 ;
            rom[27026] = 8'hec ;
            rom[27027] = 8'he6 ;
            rom[27028] = 8'h0a ;
            rom[27029] = 8'hf3 ;
            rom[27030] = 8'h1b ;
            rom[27031] = 8'hd2 ;
            rom[27032] = 8'h04 ;
            rom[27033] = 8'h17 ;
            rom[27034] = 8'h09 ;
            rom[27035] = 8'h22 ;
            rom[27036] = 8'h1e ;
            rom[27037] = 8'hff ;
            rom[27038] = 8'h10 ;
            rom[27039] = 8'hff ;
            rom[27040] = 8'h15 ;
            rom[27041] = 8'hb9 ;
            rom[27042] = 8'hd1 ;
            rom[27043] = 8'hfd ;
            rom[27044] = 8'h00 ;
            rom[27045] = 8'he1 ;
            rom[27046] = 8'hfc ;
            rom[27047] = 8'hf9 ;
            rom[27048] = 8'h0f ;
            rom[27049] = 8'h01 ;
            rom[27050] = 8'h1e ;
            rom[27051] = 8'hfe ;
            rom[27052] = 8'hfd ;
            rom[27053] = 8'hf5 ;
            rom[27054] = 8'hea ;
            rom[27055] = 8'h1d ;
            rom[27056] = 8'he0 ;
            rom[27057] = 8'h02 ;
            rom[27058] = 8'h0f ;
            rom[27059] = 8'hf8 ;
            rom[27060] = 8'hf7 ;
            rom[27061] = 8'heb ;
            rom[27062] = 8'hdd ;
            rom[27063] = 8'he0 ;
            rom[27064] = 8'hfe ;
            rom[27065] = 8'h29 ;
            rom[27066] = 8'h0a ;
            rom[27067] = 8'h23 ;
            rom[27068] = 8'hbb ;
            rom[27069] = 8'h08 ;
            rom[27070] = 8'hfc ;
            rom[27071] = 8'h19 ;
            rom[27072] = 8'hf3 ;
            rom[27073] = 8'hee ;
            rom[27074] = 8'hf7 ;
            rom[27075] = 8'he8 ;
            rom[27076] = 8'h03 ;
            rom[27077] = 8'hce ;
            rom[27078] = 8'hfc ;
            rom[27079] = 8'hd5 ;
            rom[27080] = 8'h14 ;
            rom[27081] = 8'hde ;
            rom[27082] = 8'hf9 ;
            rom[27083] = 8'h2f ;
            rom[27084] = 8'he5 ;
            rom[27085] = 8'h05 ;
            rom[27086] = 8'h06 ;
            rom[27087] = 8'h0b ;
            rom[27088] = 8'h2b ;
            rom[27089] = 8'hf8 ;
            rom[27090] = 8'hec ;
            rom[27091] = 8'hfd ;
            rom[27092] = 8'he6 ;
            rom[27093] = 8'hd9 ;
            rom[27094] = 8'h01 ;
            rom[27095] = 8'hf3 ;
            rom[27096] = 8'h05 ;
            rom[27097] = 8'hf9 ;
            rom[27098] = 8'h32 ;
            rom[27099] = 8'h16 ;
            rom[27100] = 8'h13 ;
            rom[27101] = 8'hfc ;
            rom[27102] = 8'h17 ;
            rom[27103] = 8'he7 ;
            rom[27104] = 8'hfa ;
            rom[27105] = 8'h24 ;
            rom[27106] = 8'he3 ;
            rom[27107] = 8'hd9 ;
            rom[27108] = 8'hf6 ;
            rom[27109] = 8'he7 ;
            rom[27110] = 8'hff ;
            rom[27111] = 8'h1a ;
            rom[27112] = 8'he7 ;
            rom[27113] = 8'h14 ;
            rom[27114] = 8'h01 ;
            rom[27115] = 8'hfa ;
            rom[27116] = 8'h0b ;
            rom[27117] = 8'h2c ;
            rom[27118] = 8'hf1 ;
            rom[27119] = 8'h22 ;
            rom[27120] = 8'h24 ;
            rom[27121] = 8'h21 ;
            rom[27122] = 8'h20 ;
            rom[27123] = 8'hff ;
            rom[27124] = 8'h30 ;
            rom[27125] = 8'h12 ;
            rom[27126] = 8'hf6 ;
            rom[27127] = 8'h1c ;
            rom[27128] = 8'h01 ;
            rom[27129] = 8'h12 ;
            rom[27130] = 8'h23 ;
            rom[27131] = 8'h25 ;
            rom[27132] = 8'he9 ;
            rom[27133] = 8'h20 ;
            rom[27134] = 8'h16 ;
            rom[27135] = 8'hdc ;
            rom[27136] = 8'hfd ;
            rom[27137] = 8'h0e ;
            rom[27138] = 8'hff ;
            rom[27139] = 8'h1f ;
            rom[27140] = 8'h1b ;
            rom[27141] = 8'hec ;
            rom[27142] = 8'hda ;
            rom[27143] = 8'he6 ;
            rom[27144] = 8'hfd ;
            rom[27145] = 8'hff ;
            rom[27146] = 8'hfa ;
            rom[27147] = 8'h01 ;
            rom[27148] = 8'hd3 ;
            rom[27149] = 8'hfc ;
            rom[27150] = 8'h18 ;
            rom[27151] = 8'h18 ;
            rom[27152] = 8'h03 ;
            rom[27153] = 8'h1b ;
            rom[27154] = 8'hfa ;
            rom[27155] = 8'hf4 ;
            rom[27156] = 8'h1d ;
            rom[27157] = 8'h17 ;
            rom[27158] = 8'hd4 ;
            rom[27159] = 8'h09 ;
            rom[27160] = 8'h06 ;
            rom[27161] = 8'h04 ;
            rom[27162] = 8'h1b ;
            rom[27163] = 8'hf3 ;
            rom[27164] = 8'he7 ;
            rom[27165] = 8'hdb ;
            rom[27166] = 8'hfe ;
            rom[27167] = 8'h20 ;
            rom[27168] = 8'hd4 ;
            rom[27169] = 8'h16 ;
            rom[27170] = 8'h05 ;
            rom[27171] = 8'h05 ;
            rom[27172] = 8'hf8 ;
            rom[27173] = 8'hee ;
            rom[27174] = 8'hef ;
            rom[27175] = 8'h19 ;
            rom[27176] = 8'hf0 ;
            rom[27177] = 8'h03 ;
            rom[27178] = 8'he7 ;
            rom[27179] = 8'hed ;
            rom[27180] = 8'hf2 ;
            rom[27181] = 8'hfb ;
            rom[27182] = 8'h17 ;
            rom[27183] = 8'hd9 ;
            rom[27184] = 8'h12 ;
            rom[27185] = 8'hf6 ;
            rom[27186] = 8'hca ;
            rom[27187] = 8'h08 ;
            rom[27188] = 8'h1c ;
            rom[27189] = 8'hc1 ;
            rom[27190] = 8'hf1 ;
            rom[27191] = 8'h00 ;
            rom[27192] = 8'h1e ;
            rom[27193] = 8'h02 ;
            rom[27194] = 8'hf1 ;
            rom[27195] = 8'hf4 ;
            rom[27196] = 8'h08 ;
            rom[27197] = 8'he6 ;
            rom[27198] = 8'hda ;
            rom[27199] = 8'hf7 ;
            rom[27200] = 8'he9 ;
            rom[27201] = 8'hf9 ;
            rom[27202] = 8'h0a ;
            rom[27203] = 8'hf8 ;
            rom[27204] = 8'h03 ;
            rom[27205] = 8'hee ;
            rom[27206] = 8'hed ;
            rom[27207] = 8'hf9 ;
            rom[27208] = 8'h06 ;
            rom[27209] = 8'h03 ;
            rom[27210] = 8'h0b ;
            rom[27211] = 8'h10 ;
            rom[27212] = 8'h23 ;
            rom[27213] = 8'hfd ;
            rom[27214] = 8'hcf ;
            rom[27215] = 8'h09 ;
            rom[27216] = 8'hf6 ;
            rom[27217] = 8'hfb ;
            rom[27218] = 8'he2 ;
            rom[27219] = 8'h05 ;
            rom[27220] = 8'h06 ;
            rom[27221] = 8'hfd ;
            rom[27222] = 8'hcf ;
            rom[27223] = 8'h15 ;
            rom[27224] = 8'hfd ;
            rom[27225] = 8'hec ;
            rom[27226] = 8'hf1 ;
            rom[27227] = 8'h08 ;
            rom[27228] = 8'h0b ;
            rom[27229] = 8'h1f ;
            rom[27230] = 8'h0c ;
            rom[27231] = 8'h26 ;
            rom[27232] = 8'hff ;
            rom[27233] = 8'ha3 ;
            rom[27234] = 8'h00 ;
            rom[27235] = 8'hfa ;
            rom[27236] = 8'hfd ;
            rom[27237] = 8'he4 ;
            rom[27238] = 8'hec ;
            rom[27239] = 8'h04 ;
            rom[27240] = 8'h91 ;
            rom[27241] = 8'hc1 ;
            rom[27242] = 8'he8 ;
            rom[27243] = 8'hec ;
            rom[27244] = 8'heb ;
            rom[27245] = 8'hd8 ;
            rom[27246] = 8'hfd ;
            rom[27247] = 8'h2e ;
            rom[27248] = 8'h1f ;
            rom[27249] = 8'he2 ;
            rom[27250] = 8'h26 ;
            rom[27251] = 8'hea ;
            rom[27252] = 8'h09 ;
            rom[27253] = 8'hfc ;
            rom[27254] = 8'hec ;
            rom[27255] = 8'hf1 ;
            rom[27256] = 8'h0b ;
            rom[27257] = 8'hf7 ;
            rom[27258] = 8'h02 ;
            rom[27259] = 8'he8 ;
            rom[27260] = 8'h09 ;
            rom[27261] = 8'hf5 ;
            rom[27262] = 8'hd4 ;
            rom[27263] = 8'hdb ;
            rom[27264] = 8'he9 ;
            rom[27265] = 8'h0a ;
            rom[27266] = 8'h16 ;
            rom[27267] = 8'hf0 ;
            rom[27268] = 8'hf4 ;
            rom[27269] = 8'hea ;
            rom[27270] = 8'h09 ;
            rom[27271] = 8'h06 ;
            rom[27272] = 8'h0e ;
            rom[27273] = 8'h0e ;
            rom[27274] = 8'hff ;
            rom[27275] = 8'h0a ;
            rom[27276] = 8'h0b ;
            rom[27277] = 8'h1b ;
            rom[27278] = 8'h1a ;
            rom[27279] = 8'hf3 ;
            rom[27280] = 8'hef ;
            rom[27281] = 8'h07 ;
            rom[27282] = 8'h10 ;
            rom[27283] = 8'hf0 ;
            rom[27284] = 8'h10 ;
            rom[27285] = 8'hdf ;
            rom[27286] = 8'h03 ;
            rom[27287] = 8'hf2 ;
            rom[27288] = 8'hfb ;
            rom[27289] = 8'hfb ;
            rom[27290] = 8'h09 ;
            rom[27291] = 8'hdf ;
            rom[27292] = 8'hf2 ;
            rom[27293] = 8'h05 ;
            rom[27294] = 8'hfa ;
            rom[27295] = 8'h0e ;
            rom[27296] = 8'hfd ;
            rom[27297] = 8'hce ;
            rom[27298] = 8'hfa ;
            rom[27299] = 8'h1a ;
            rom[27300] = 8'hf9 ;
            rom[27301] = 8'hf3 ;
            rom[27302] = 8'h11 ;
            rom[27303] = 8'hff ;
            rom[27304] = 8'hf2 ;
            rom[27305] = 8'he9 ;
            rom[27306] = 8'hdd ;
            rom[27307] = 8'h00 ;
            rom[27308] = 8'he0 ;
            rom[27309] = 8'h0f ;
            rom[27310] = 8'hfc ;
            rom[27311] = 8'h07 ;
            rom[27312] = 8'h02 ;
            rom[27313] = 8'h14 ;
            rom[27314] = 8'h1c ;
            rom[27315] = 8'hf6 ;
            rom[27316] = 8'h09 ;
            rom[27317] = 8'h1a ;
            rom[27318] = 8'hfd ;
            rom[27319] = 8'hbc ;
            rom[27320] = 8'h04 ;
            rom[27321] = 8'h05 ;
            rom[27322] = 8'h00 ;
            rom[27323] = 8'h0f ;
            rom[27324] = 8'he9 ;
            rom[27325] = 8'hf9 ;
            rom[27326] = 8'hff ;
            rom[27327] = 8'he3 ;
            rom[27328] = 8'h1d ;
            rom[27329] = 8'heb ;
            rom[27330] = 8'h07 ;
            rom[27331] = 8'hf9 ;
            rom[27332] = 8'hee ;
            rom[27333] = 8'h11 ;
            rom[27334] = 8'hd0 ;
            rom[27335] = 8'he5 ;
            rom[27336] = 8'he5 ;
            rom[27337] = 8'hf2 ;
            rom[27338] = 8'hf7 ;
            rom[27339] = 8'h09 ;
            rom[27340] = 8'h09 ;
            rom[27341] = 8'hf4 ;
            rom[27342] = 8'hec ;
            rom[27343] = 8'hf7 ;
            rom[27344] = 8'hd9 ;
            rom[27345] = 8'hf8 ;
            rom[27346] = 8'h0d ;
            rom[27347] = 8'hdf ;
            rom[27348] = 8'heb ;
            rom[27349] = 8'h02 ;
            rom[27350] = 8'h0d ;
            rom[27351] = 8'hec ;
            rom[27352] = 8'hfb ;
            rom[27353] = 8'hf1 ;
            rom[27354] = 8'hf4 ;
            rom[27355] = 8'h0d ;
            rom[27356] = 8'hee ;
            rom[27357] = 8'h17 ;
            rom[27358] = 8'he2 ;
            rom[27359] = 8'hdb ;
            rom[27360] = 8'h03 ;
            rom[27361] = 8'hfa ;
            rom[27362] = 8'he6 ;
            rom[27363] = 8'h04 ;
            rom[27364] = 8'h1c ;
            rom[27365] = 8'h11 ;
            rom[27366] = 8'hdc ;
            rom[27367] = 8'ha8 ;
            rom[27368] = 8'h25 ;
            rom[27369] = 8'h09 ;
            rom[27370] = 8'hfe ;
            rom[27371] = 8'h0a ;
            rom[27372] = 8'hb2 ;
            rom[27373] = 8'h04 ;
            rom[27374] = 8'hfe ;
            rom[27375] = 8'h14 ;
            rom[27376] = 8'he9 ;
            rom[27377] = 8'hf9 ;
            rom[27378] = 8'h01 ;
            rom[27379] = 8'hf9 ;
            rom[27380] = 8'h02 ;
            rom[27381] = 8'hda ;
            rom[27382] = 8'h07 ;
            rom[27383] = 8'hf0 ;
            rom[27384] = 8'hd7 ;
            rom[27385] = 8'h08 ;
            rom[27386] = 8'h12 ;
            rom[27387] = 8'h02 ;
            rom[27388] = 8'hd9 ;
            rom[27389] = 8'hcb ;
            rom[27390] = 8'hd3 ;
            rom[27391] = 8'hf2 ;
            rom[27392] = 8'h16 ;
            rom[27393] = 8'h0e ;
            rom[27394] = 8'hef ;
            rom[27395] = 8'he7 ;
            rom[27396] = 8'hf9 ;
            rom[27397] = 8'hd2 ;
            rom[27398] = 8'hc0 ;
            rom[27399] = 8'h0a ;
            rom[27400] = 8'h10 ;
            rom[27401] = 8'hf8 ;
            rom[27402] = 8'hfe ;
            rom[27403] = 8'hf5 ;
            rom[27404] = 8'hba ;
            rom[27405] = 8'h09 ;
            rom[27406] = 8'h18 ;
            rom[27407] = 8'h0b ;
            rom[27408] = 8'h0f ;
            rom[27409] = 8'hf9 ;
            rom[27410] = 8'hf8 ;
            rom[27411] = 8'h1d ;
            rom[27412] = 8'hd6 ;
            rom[27413] = 8'h0c ;
            rom[27414] = 8'h08 ;
            rom[27415] = 8'h11 ;
            rom[27416] = 8'hf7 ;
            rom[27417] = 8'h04 ;
            rom[27418] = 8'hee ;
            rom[27419] = 8'hf8 ;
            rom[27420] = 8'h19 ;
            rom[27421] = 8'h1e ;
            rom[27422] = 8'h17 ;
            rom[27423] = 8'hdc ;
            rom[27424] = 8'hcd ;
            rom[27425] = 8'h1f ;
            rom[27426] = 8'h0a ;
            rom[27427] = 8'hff ;
            rom[27428] = 8'h05 ;
            rom[27429] = 8'he8 ;
            rom[27430] = 8'hbe ;
            rom[27431] = 8'h0d ;
            rom[27432] = 8'hfc ;
            rom[27433] = 8'h0b ;
            rom[27434] = 8'hf9 ;
            rom[27435] = 8'hf9 ;
            rom[27436] = 8'hd9 ;
            rom[27437] = 8'hed ;
            rom[27438] = 8'he0 ;
            rom[27439] = 8'h02 ;
            rom[27440] = 8'h16 ;
            rom[27441] = 8'h0d ;
            rom[27442] = 8'hed ;
            rom[27443] = 8'hce ;
            rom[27444] = 8'hdf ;
            rom[27445] = 8'hfd ;
            rom[27446] = 8'h0d ;
            rom[27447] = 8'he7 ;
            rom[27448] = 8'h27 ;
            rom[27449] = 8'h0c ;
            rom[27450] = 8'h03 ;
            rom[27451] = 8'h05 ;
            rom[27452] = 8'h09 ;
            rom[27453] = 8'hf0 ;
            rom[27454] = 8'hfb ;
            rom[27455] = 8'hc6 ;
            rom[27456] = 8'hc3 ;
            rom[27457] = 8'he2 ;
            rom[27458] = 8'he5 ;
            rom[27459] = 8'hf3 ;
            rom[27460] = 8'h05 ;
            rom[27461] = 8'h0b ;
            rom[27462] = 8'hf4 ;
            rom[27463] = 8'he3 ;
            rom[27464] = 8'h06 ;
            rom[27465] = 8'h06 ;
            rom[27466] = 8'hea ;
            rom[27467] = 8'hd0 ;
            rom[27468] = 8'hf5 ;
            rom[27469] = 8'h1f ;
            rom[27470] = 8'hee ;
            rom[27471] = 8'hc6 ;
            rom[27472] = 8'heb ;
            rom[27473] = 8'hee ;
            rom[27474] = 8'hff ;
            rom[27475] = 8'hf7 ;
            rom[27476] = 8'hfc ;
            rom[27477] = 8'he6 ;
            rom[27478] = 8'h13 ;
            rom[27479] = 8'h0c ;
            rom[27480] = 8'hf8 ;
            rom[27481] = 8'hf8 ;
            rom[27482] = 8'he1 ;
            rom[27483] = 8'h00 ;
            rom[27484] = 8'h08 ;
            rom[27485] = 8'h05 ;
            rom[27486] = 8'he7 ;
            rom[27487] = 8'he1 ;
            rom[27488] = 8'hfe ;
            rom[27489] = 8'hee ;
            rom[27490] = 8'hf4 ;
            rom[27491] = 8'h0d ;
            rom[27492] = 8'h0d ;
            rom[27493] = 8'h07 ;
            rom[27494] = 8'hec ;
            rom[27495] = 8'hee ;
            rom[27496] = 8'hcc ;
            rom[27497] = 8'h0c ;
            rom[27498] = 8'hf9 ;
            rom[27499] = 8'hea ;
            rom[27500] = 8'hfe ;
            rom[27501] = 8'h1b ;
            rom[27502] = 8'he7 ;
            rom[27503] = 8'hdc ;
            rom[27504] = 8'hd3 ;
            rom[27505] = 8'hdf ;
            rom[27506] = 8'he5 ;
            rom[27507] = 8'hfb ;
            rom[27508] = 8'he3 ;
            rom[27509] = 8'h18 ;
            rom[27510] = 8'he9 ;
            rom[27511] = 8'hda ;
            rom[27512] = 8'h04 ;
            rom[27513] = 8'hfb ;
            rom[27514] = 8'hca ;
            rom[27515] = 8'h18 ;
            rom[27516] = 8'h04 ;
            rom[27517] = 8'hff ;
            rom[27518] = 8'h2a ;
            rom[27519] = 8'hdf ;
            rom[27520] = 8'h38 ;
            rom[27521] = 8'he5 ;
            rom[27522] = 8'he6 ;
            rom[27523] = 8'h28 ;
            rom[27524] = 8'hf3 ;
            rom[27525] = 8'he8 ;
            rom[27526] = 8'hf9 ;
            rom[27527] = 8'h0d ;
            rom[27528] = 8'he9 ;
            rom[27529] = 8'h1a ;
            rom[27530] = 8'hce ;
            rom[27531] = 8'h15 ;
            rom[27532] = 8'h0c ;
            rom[27533] = 8'h0c ;
            rom[27534] = 8'hcb ;
            rom[27535] = 8'h13 ;
            rom[27536] = 8'h02 ;
            rom[27537] = 8'h19 ;
            rom[27538] = 8'h22 ;
            rom[27539] = 8'h06 ;
            rom[27540] = 8'h11 ;
            rom[27541] = 8'hdb ;
            rom[27542] = 8'h04 ;
            rom[27543] = 8'h0d ;
            rom[27544] = 8'h04 ;
            rom[27545] = 8'h18 ;
            rom[27546] = 8'he0 ;
            rom[27547] = 8'h13 ;
            rom[27548] = 8'hf3 ;
            rom[27549] = 8'h06 ;
            rom[27550] = 8'h03 ;
            rom[27551] = 8'hff ;
            rom[27552] = 8'hc7 ;
            rom[27553] = 8'hde ;
            rom[27554] = 8'hfc ;
            rom[27555] = 8'hf5 ;
            rom[27556] = 8'hcc ;
            rom[27557] = 8'hfd ;
            rom[27558] = 8'hf8 ;
            rom[27559] = 8'he4 ;
            rom[27560] = 8'hf4 ;
            rom[27561] = 8'hf5 ;
            rom[27562] = 8'hf9 ;
            rom[27563] = 8'ha8 ;
            rom[27564] = 8'h17 ;
            rom[27565] = 8'h13 ;
            rom[27566] = 8'hf0 ;
            rom[27567] = 8'h10 ;
            rom[27568] = 8'h15 ;
            rom[27569] = 8'heb ;
            rom[27570] = 8'h08 ;
            rom[27571] = 8'h1d ;
            rom[27572] = 8'hf7 ;
            rom[27573] = 8'he1 ;
            rom[27574] = 8'h07 ;
            rom[27575] = 8'he0 ;
            rom[27576] = 8'h12 ;
            rom[27577] = 8'h16 ;
            rom[27578] = 8'hf3 ;
            rom[27579] = 8'h10 ;
            rom[27580] = 8'hcc ;
            rom[27581] = 8'h08 ;
            rom[27582] = 8'he7 ;
            rom[27583] = 8'h1b ;
            rom[27584] = 8'hdf ;
            rom[27585] = 8'hf1 ;
            rom[27586] = 8'hf4 ;
            rom[27587] = 8'h07 ;
            rom[27588] = 8'he5 ;
            rom[27589] = 8'hf2 ;
            rom[27590] = 8'hef ;
            rom[27591] = 8'hd2 ;
            rom[27592] = 8'hd0 ;
            rom[27593] = 8'hf7 ;
            rom[27594] = 8'h3b ;
            rom[27595] = 8'h0f ;
            rom[27596] = 8'h16 ;
            rom[27597] = 8'h17 ;
            rom[27598] = 8'h12 ;
            rom[27599] = 8'h04 ;
            rom[27600] = 8'h02 ;
            rom[27601] = 8'h18 ;
            rom[27602] = 8'hd8 ;
            rom[27603] = 8'hef ;
            rom[27604] = 8'hf3 ;
            rom[27605] = 8'hf4 ;
            rom[27606] = 8'hd2 ;
            rom[27607] = 8'hf7 ;
            rom[27608] = 8'h0a ;
            rom[27609] = 8'hfd ;
            rom[27610] = 8'hea ;
            rom[27611] = 8'h1b ;
            rom[27612] = 8'h20 ;
            rom[27613] = 8'hda ;
            rom[27614] = 8'h09 ;
            rom[27615] = 8'h05 ;
            rom[27616] = 8'h1a ;
            rom[27617] = 8'h0a ;
            rom[27618] = 8'hf9 ;
            rom[27619] = 8'hf0 ;
            rom[27620] = 8'h0c ;
            rom[27621] = 8'h06 ;
            rom[27622] = 8'hda ;
            rom[27623] = 8'hf0 ;
            rom[27624] = 8'h0e ;
            rom[27625] = 8'h06 ;
            rom[27626] = 8'hee ;
            rom[27627] = 8'h0f ;
            rom[27628] = 8'hed ;
            rom[27629] = 8'h00 ;
            rom[27630] = 8'hbe ;
            rom[27631] = 8'he3 ;
            rom[27632] = 8'h06 ;
            rom[27633] = 8'hff ;
            rom[27634] = 8'hfd ;
            rom[27635] = 8'he2 ;
            rom[27636] = 8'h0b ;
            rom[27637] = 8'hf1 ;
            rom[27638] = 8'h02 ;
            rom[27639] = 8'h19 ;
            rom[27640] = 8'h08 ;
            rom[27641] = 8'hd7 ;
            rom[27642] = 8'hf3 ;
            rom[27643] = 8'h23 ;
            rom[27644] = 8'h03 ;
            rom[27645] = 8'hea ;
            rom[27646] = 8'hf4 ;
            rom[27647] = 8'hfb ;
            rom[27648] = 8'hd3 ;
            rom[27649] = 8'h03 ;
            rom[27650] = 8'hf6 ;
            rom[27651] = 8'h06 ;
            rom[27652] = 8'hfb ;
            rom[27653] = 8'hf8 ;
            rom[27654] = 8'h0a ;
            rom[27655] = 8'h1d ;
            rom[27656] = 8'h03 ;
            rom[27657] = 8'h16 ;
            rom[27658] = 8'h00 ;
            rom[27659] = 8'h1a ;
            rom[27660] = 8'h15 ;
            rom[27661] = 8'he8 ;
            rom[27662] = 8'he8 ;
            rom[27663] = 8'h07 ;
            rom[27664] = 8'h11 ;
            rom[27665] = 8'hdb ;
            rom[27666] = 8'h0b ;
            rom[27667] = 8'h0a ;
            rom[27668] = 8'h16 ;
            rom[27669] = 8'hf3 ;
            rom[27670] = 8'h06 ;
            rom[27671] = 8'h0d ;
            rom[27672] = 8'h15 ;
            rom[27673] = 8'hf6 ;
            rom[27674] = 8'hf4 ;
            rom[27675] = 8'hf7 ;
            rom[27676] = 8'hfb ;
            rom[27677] = 8'hde ;
            rom[27678] = 8'hec ;
            rom[27679] = 8'hf6 ;
            rom[27680] = 8'h05 ;
            rom[27681] = 8'h01 ;
            rom[27682] = 8'hfd ;
            rom[27683] = 8'h07 ;
            rom[27684] = 8'hfe ;
            rom[27685] = 8'h07 ;
            rom[27686] = 8'hdb ;
            rom[27687] = 8'heb ;
            rom[27688] = 8'h0c ;
            rom[27689] = 8'hdc ;
            rom[27690] = 8'h08 ;
            rom[27691] = 8'hf7 ;
            rom[27692] = 8'h18 ;
            rom[27693] = 8'h22 ;
            rom[27694] = 8'hdf ;
            rom[27695] = 8'he7 ;
            rom[27696] = 8'h03 ;
            rom[27697] = 8'h06 ;
            rom[27698] = 8'h0e ;
            rom[27699] = 8'h00 ;
            rom[27700] = 8'hf5 ;
            rom[27701] = 8'hf5 ;
            rom[27702] = 8'h01 ;
            rom[27703] = 8'hcf ;
            rom[27704] = 8'h1b ;
            rom[27705] = 8'h2b ;
            rom[27706] = 8'h04 ;
            rom[27707] = 8'h11 ;
            rom[27708] = 8'h02 ;
            rom[27709] = 8'h31 ;
            rom[27710] = 8'h03 ;
            rom[27711] = 8'h0f ;
            rom[27712] = 8'h1a ;
            rom[27713] = 8'hed ;
            rom[27714] = 8'hf2 ;
            rom[27715] = 8'hdf ;
            rom[27716] = 8'hf1 ;
            rom[27717] = 8'h06 ;
            rom[27718] = 8'hd5 ;
            rom[27719] = 8'hee ;
            rom[27720] = 8'he5 ;
            rom[27721] = 8'h01 ;
            rom[27722] = 8'hf0 ;
            rom[27723] = 8'hf5 ;
            rom[27724] = 8'hff ;
            rom[27725] = 8'h15 ;
            rom[27726] = 8'h02 ;
            rom[27727] = 8'h1a ;
            rom[27728] = 8'h24 ;
            rom[27729] = 8'hfd ;
            rom[27730] = 8'hf5 ;
            rom[27731] = 8'hdd ;
            rom[27732] = 8'hef ;
            rom[27733] = 8'ha9 ;
            rom[27734] = 8'hfa ;
            rom[27735] = 8'hbd ;
            rom[27736] = 8'h15 ;
            rom[27737] = 8'h14 ;
            rom[27738] = 8'h34 ;
            rom[27739] = 8'heb ;
            rom[27740] = 8'hea ;
            rom[27741] = 8'h04 ;
            rom[27742] = 8'h02 ;
            rom[27743] = 8'h07 ;
            rom[27744] = 8'h1b ;
            rom[27745] = 8'h04 ;
            rom[27746] = 8'h14 ;
            rom[27747] = 8'h1e ;
            rom[27748] = 8'h26 ;
            rom[27749] = 8'hec ;
            rom[27750] = 8'hff ;
            rom[27751] = 8'h08 ;
            rom[27752] = 8'h03 ;
            rom[27753] = 8'hff ;
            rom[27754] = 8'hf3 ;
            rom[27755] = 8'h1e ;
            rom[27756] = 8'he9 ;
            rom[27757] = 8'h31 ;
            rom[27758] = 8'hf6 ;
            rom[27759] = 8'hed ;
            rom[27760] = 8'hfa ;
            rom[27761] = 8'h0d ;
            rom[27762] = 8'hee ;
            rom[27763] = 8'hf5 ;
            rom[27764] = 8'h17 ;
            rom[27765] = 8'hef ;
            rom[27766] = 8'h0f ;
            rom[27767] = 8'h3e ;
            rom[27768] = 8'h10 ;
            rom[27769] = 8'hfa ;
            rom[27770] = 8'hf7 ;
            rom[27771] = 8'hd5 ;
            rom[27772] = 8'he5 ;
            rom[27773] = 8'he8 ;
            rom[27774] = 8'he0 ;
            rom[27775] = 8'h14 ;
            rom[27776] = 8'h13 ;
            rom[27777] = 8'h21 ;
            rom[27778] = 8'hfc ;
            rom[27779] = 8'hd5 ;
            rom[27780] = 8'h1f ;
            rom[27781] = 8'hff ;
            rom[27782] = 8'hdd ;
            rom[27783] = 8'h12 ;
            rom[27784] = 8'hfa ;
            rom[27785] = 8'hf5 ;
            rom[27786] = 8'hfc ;
            rom[27787] = 8'hfe ;
            rom[27788] = 8'hf5 ;
            rom[27789] = 8'hce ;
            rom[27790] = 8'hf4 ;
            rom[27791] = 8'hf6 ;
            rom[27792] = 8'h08 ;
            rom[27793] = 8'h01 ;
            rom[27794] = 8'h04 ;
            rom[27795] = 8'h07 ;
            rom[27796] = 8'h1a ;
            rom[27797] = 8'h17 ;
            rom[27798] = 8'h21 ;
            rom[27799] = 8'he2 ;
            rom[27800] = 8'hde ;
            rom[27801] = 8'hec ;
            rom[27802] = 8'h00 ;
            rom[27803] = 8'h09 ;
            rom[27804] = 8'h22 ;
            rom[27805] = 8'h0e ;
            rom[27806] = 8'h12 ;
            rom[27807] = 8'hf1 ;
            rom[27808] = 8'h03 ;
            rom[27809] = 8'h16 ;
            rom[27810] = 8'h13 ;
            rom[27811] = 8'h20 ;
            rom[27812] = 8'h1a ;
            rom[27813] = 8'hfb ;
            rom[27814] = 8'hca ;
            rom[27815] = 8'hfb ;
            rom[27816] = 8'hf5 ;
            rom[27817] = 8'hc8 ;
            rom[27818] = 8'hfc ;
            rom[27819] = 8'h09 ;
            rom[27820] = 8'hea ;
            rom[27821] = 8'ha0 ;
            rom[27822] = 8'he2 ;
            rom[27823] = 8'h0d ;
            rom[27824] = 8'h17 ;
            rom[27825] = 8'hf5 ;
            rom[27826] = 8'h0c ;
            rom[27827] = 8'hfb ;
            rom[27828] = 8'hc2 ;
            rom[27829] = 8'h04 ;
            rom[27830] = 8'h15 ;
            rom[27831] = 8'he3 ;
            rom[27832] = 8'hed ;
            rom[27833] = 8'hf9 ;
            rom[27834] = 8'hf1 ;
            rom[27835] = 8'h07 ;
            rom[27836] = 8'h16 ;
            rom[27837] = 8'hf3 ;
            rom[27838] = 8'hf7 ;
            rom[27839] = 8'hed ;
            rom[27840] = 8'he2 ;
            rom[27841] = 8'hf6 ;
            rom[27842] = 8'hfa ;
            rom[27843] = 8'h22 ;
            rom[27844] = 8'hc6 ;
            rom[27845] = 8'hf5 ;
            rom[27846] = 8'hf5 ;
            rom[27847] = 8'h11 ;
            rom[27848] = 8'hfa ;
            rom[27849] = 8'h0c ;
            rom[27850] = 8'he9 ;
            rom[27851] = 8'h0c ;
            rom[27852] = 8'h03 ;
            rom[27853] = 8'he6 ;
            rom[27854] = 8'h06 ;
            rom[27855] = 8'he0 ;
            rom[27856] = 8'h05 ;
            rom[27857] = 8'h0c ;
            rom[27858] = 8'h05 ;
            rom[27859] = 8'hb8 ;
            rom[27860] = 8'h1f ;
            rom[27861] = 8'hca ;
            rom[27862] = 8'h09 ;
            rom[27863] = 8'hda ;
            rom[27864] = 8'h0a ;
            rom[27865] = 8'h10 ;
            rom[27866] = 8'h13 ;
            rom[27867] = 8'hf0 ;
            rom[27868] = 8'hf7 ;
            rom[27869] = 8'hec ;
            rom[27870] = 8'he7 ;
            rom[27871] = 8'he3 ;
            rom[27872] = 8'h0a ;
            rom[27873] = 8'h01 ;
            rom[27874] = 8'h01 ;
            rom[27875] = 8'he4 ;
            rom[27876] = 8'h03 ;
            rom[27877] = 8'hf1 ;
            rom[27878] = 8'hfe ;
            rom[27879] = 8'h15 ;
            rom[27880] = 8'hf1 ;
            rom[27881] = 8'h07 ;
            rom[27882] = 8'he8 ;
            rom[27883] = 8'h0e ;
            rom[27884] = 8'hdb ;
            rom[27885] = 8'h0b ;
            rom[27886] = 8'hfb ;
            rom[27887] = 8'hb8 ;
            rom[27888] = 8'h05 ;
            rom[27889] = 8'hf2 ;
            rom[27890] = 8'hf0 ;
            rom[27891] = 8'h0f ;
            rom[27892] = 8'he2 ;
            rom[27893] = 8'hf7 ;
            rom[27894] = 8'h17 ;
            rom[27895] = 8'hfe ;
            rom[27896] = 8'h0b ;
            rom[27897] = 8'hf2 ;
            rom[27898] = 8'hdc ;
            rom[27899] = 8'h2e ;
            rom[27900] = 8'he8 ;
            rom[27901] = 8'heb ;
            rom[27902] = 8'h10 ;
            rom[27903] = 8'hf0 ;
            rom[27904] = 8'h19 ;
            rom[27905] = 8'hf2 ;
            rom[27906] = 8'h08 ;
            rom[27907] = 8'h00 ;
            rom[27908] = 8'hf5 ;
            rom[27909] = 8'h06 ;
            rom[27910] = 8'h39 ;
            rom[27911] = 8'h0b ;
            rom[27912] = 8'he8 ;
            rom[27913] = 8'h26 ;
            rom[27914] = 8'hf9 ;
            rom[27915] = 8'h0e ;
            rom[27916] = 8'h01 ;
            rom[27917] = 8'h1a ;
            rom[27918] = 8'hf2 ;
            rom[27919] = 8'h06 ;
            rom[27920] = 8'he5 ;
            rom[27921] = 8'h09 ;
            rom[27922] = 8'h0d ;
            rom[27923] = 8'hec ;
            rom[27924] = 8'h04 ;
            rom[27925] = 8'h07 ;
            rom[27926] = 8'h0c ;
            rom[27927] = 8'hf8 ;
            rom[27928] = 8'he5 ;
            rom[27929] = 8'hf5 ;
            rom[27930] = 8'hf8 ;
            rom[27931] = 8'hd6 ;
            rom[27932] = 8'hf5 ;
            rom[27933] = 8'h01 ;
            rom[27934] = 8'heb ;
            rom[27935] = 8'h07 ;
            rom[27936] = 8'h28 ;
            rom[27937] = 8'h25 ;
            rom[27938] = 8'h05 ;
            rom[27939] = 8'h20 ;
            rom[27940] = 8'h1e ;
            rom[27941] = 8'hf4 ;
            rom[27942] = 8'h07 ;
            rom[27943] = 8'he8 ;
            rom[27944] = 8'hf1 ;
            rom[27945] = 8'hfa ;
            rom[27946] = 8'hce ;
            rom[27947] = 8'hf9 ;
            rom[27948] = 8'h14 ;
            rom[27949] = 8'h12 ;
            rom[27950] = 8'hf7 ;
            rom[27951] = 8'h06 ;
            rom[27952] = 8'hf6 ;
            rom[27953] = 8'hd0 ;
            rom[27954] = 8'h22 ;
            rom[27955] = 8'h00 ;
            rom[27956] = 8'hed ;
            rom[27957] = 8'hfd ;
            rom[27958] = 8'h0a ;
            rom[27959] = 8'h00 ;
            rom[27960] = 8'hfd ;
            rom[27961] = 8'hf5 ;
            rom[27962] = 8'hf9 ;
            rom[27963] = 8'h21 ;
            rom[27964] = 8'hf2 ;
            rom[27965] = 8'h0d ;
            rom[27966] = 8'h1d ;
            rom[27967] = 8'h07 ;
            rom[27968] = 8'h00 ;
            rom[27969] = 8'hfd ;
            rom[27970] = 8'h24 ;
            rom[27971] = 8'hcd ;
            rom[27972] = 8'he9 ;
            rom[27973] = 8'hfa ;
            rom[27974] = 8'he9 ;
            rom[27975] = 8'h08 ;
            rom[27976] = 8'hfc ;
            rom[27977] = 8'h24 ;
            rom[27978] = 8'h0a ;
            rom[27979] = 8'hf4 ;
            rom[27980] = 8'h08 ;
            rom[27981] = 8'h07 ;
            rom[27982] = 8'hf9 ;
            rom[27983] = 8'h18 ;
            rom[27984] = 8'hfb ;
            rom[27985] = 8'h1c ;
            rom[27986] = 8'hed ;
            rom[27987] = 8'hfd ;
            rom[27988] = 8'h10 ;
            rom[27989] = 8'h1d ;
            rom[27990] = 8'hcd ;
            rom[27991] = 8'h05 ;
            rom[27992] = 8'hf1 ;
            rom[27993] = 8'hfa ;
            rom[27994] = 8'h1b ;
            rom[27995] = 8'h00 ;
            rom[27996] = 8'hf1 ;
            rom[27997] = 8'he8 ;
            rom[27998] = 8'h09 ;
            rom[27999] = 8'h0b ;
            rom[28000] = 8'hfb ;
            rom[28001] = 8'hdf ;
            rom[28002] = 8'h26 ;
            rom[28003] = 8'h15 ;
            rom[28004] = 8'h15 ;
            rom[28005] = 8'hf2 ;
            rom[28006] = 8'hfc ;
            rom[28007] = 8'hfe ;
            rom[28008] = 8'h16 ;
            rom[28009] = 8'h01 ;
            rom[28010] = 8'h04 ;
            rom[28011] = 8'h21 ;
            rom[28012] = 8'hf8 ;
            rom[28013] = 8'hff ;
            rom[28014] = 8'h2d ;
            rom[28015] = 8'h19 ;
            rom[28016] = 8'h00 ;
            rom[28017] = 8'hf0 ;
            rom[28018] = 8'hcd ;
            rom[28019] = 8'h15 ;
            rom[28020] = 8'h35 ;
            rom[28021] = 8'heb ;
            rom[28022] = 8'h1e ;
            rom[28023] = 8'h22 ;
            rom[28024] = 8'h04 ;
            rom[28025] = 8'h18 ;
            rom[28026] = 8'h0f ;
            rom[28027] = 8'h10 ;
            rom[28028] = 8'h12 ;
            rom[28029] = 8'hf8 ;
            rom[28030] = 8'hf1 ;
            rom[28031] = 8'h18 ;
            rom[28032] = 8'h0e ;
            rom[28033] = 8'hf2 ;
            rom[28034] = 8'hf6 ;
            rom[28035] = 8'h20 ;
            rom[28036] = 8'h0a ;
            rom[28037] = 8'hd4 ;
            rom[28038] = 8'hf4 ;
            rom[28039] = 8'h21 ;
            rom[28040] = 8'hfe ;
            rom[28041] = 8'h0b ;
            rom[28042] = 8'h1c ;
            rom[28043] = 8'hbf ;
            rom[28044] = 8'hdb ;
            rom[28045] = 8'hd6 ;
            rom[28046] = 8'h22 ;
            rom[28047] = 8'hea ;
            rom[28048] = 8'hf8 ;
            rom[28049] = 8'hff ;
            rom[28050] = 8'h0b ;
            rom[28051] = 8'hd3 ;
            rom[28052] = 8'hea ;
            rom[28053] = 8'hd3 ;
            rom[28054] = 8'hfd ;
            rom[28055] = 8'hc8 ;
            rom[28056] = 8'hef ;
            rom[28057] = 8'hf0 ;
            rom[28058] = 8'hfc ;
            rom[28059] = 8'h04 ;
            rom[28060] = 8'h1c ;
            rom[28061] = 8'h0a ;
            rom[28062] = 8'hf6 ;
            rom[28063] = 8'h07 ;
            rom[28064] = 8'hf6 ;
            rom[28065] = 8'hf5 ;
            rom[28066] = 8'hf4 ;
            rom[28067] = 8'h0e ;
            rom[28068] = 8'hec ;
            rom[28069] = 8'h16 ;
            rom[28070] = 8'he7 ;
            rom[28071] = 8'h21 ;
            rom[28072] = 8'hc8 ;
            rom[28073] = 8'h1c ;
            rom[28074] = 8'hf8 ;
            rom[28075] = 8'h0e ;
            rom[28076] = 8'h01 ;
            rom[28077] = 8'hdb ;
            rom[28078] = 8'hdb ;
            rom[28079] = 8'h13 ;
            rom[28080] = 8'h1e ;
            rom[28081] = 8'h02 ;
            rom[28082] = 8'hff ;
            rom[28083] = 8'hff ;
            rom[28084] = 8'he0 ;
            rom[28085] = 8'hfa ;
            rom[28086] = 8'hff ;
            rom[28087] = 8'h12 ;
            rom[28088] = 8'h0a ;
            rom[28089] = 8'hed ;
            rom[28090] = 8'h08 ;
            rom[28091] = 8'h16 ;
            rom[28092] = 8'hf9 ;
            rom[28093] = 8'hf9 ;
            rom[28094] = 8'h0b ;
            rom[28095] = 8'hfd ;
            rom[28096] = 8'h0b ;
            rom[28097] = 8'h00 ;
            rom[28098] = 8'hdb ;
            rom[28099] = 8'he4 ;
            rom[28100] = 8'hf5 ;
            rom[28101] = 8'hed ;
            rom[28102] = 8'hfa ;
            rom[28103] = 8'hc5 ;
            rom[28104] = 8'h17 ;
            rom[28105] = 8'hf9 ;
            rom[28106] = 8'hf7 ;
            rom[28107] = 8'hf3 ;
            rom[28108] = 8'hf8 ;
            rom[28109] = 8'hfc ;
            rom[28110] = 8'he4 ;
            rom[28111] = 8'hd9 ;
            rom[28112] = 8'h00 ;
            rom[28113] = 8'hbd ;
            rom[28114] = 8'h0b ;
            rom[28115] = 8'hcd ;
            rom[28116] = 8'hfa ;
            rom[28117] = 8'h06 ;
            rom[28118] = 8'he8 ;
            rom[28119] = 8'hff ;
            rom[28120] = 8'h1f ;
            rom[28121] = 8'h05 ;
            rom[28122] = 8'h01 ;
            rom[28123] = 8'h17 ;
            rom[28124] = 8'h18 ;
            rom[28125] = 8'hd3 ;
            rom[28126] = 8'hbb ;
            rom[28127] = 8'h16 ;
            rom[28128] = 8'hf9 ;
            rom[28129] = 8'h19 ;
            rom[28130] = 8'h1f ;
            rom[28131] = 8'hfc ;
            rom[28132] = 8'he6 ;
            rom[28133] = 8'h05 ;
            rom[28134] = 8'h00 ;
            rom[28135] = 8'hf3 ;
            rom[28136] = 8'hbf ;
            rom[28137] = 8'hf4 ;
            rom[28138] = 8'hf0 ;
            rom[28139] = 8'hfc ;
            rom[28140] = 8'hf4 ;
            rom[28141] = 8'hfd ;
            rom[28142] = 8'he6 ;
            rom[28143] = 8'hff ;
            rom[28144] = 8'hf9 ;
            rom[28145] = 8'hdf ;
            rom[28146] = 8'hf3 ;
            rom[28147] = 8'h0a ;
            rom[28148] = 8'he9 ;
            rom[28149] = 8'h18 ;
            rom[28150] = 8'he0 ;
            rom[28151] = 8'h09 ;
            rom[28152] = 8'hf7 ;
            rom[28153] = 8'h0f ;
            rom[28154] = 8'hc4 ;
            rom[28155] = 8'h17 ;
            rom[28156] = 8'hfe ;
            rom[28157] = 8'h16 ;
            rom[28158] = 8'h06 ;
            rom[28159] = 8'h19 ;
            rom[28160] = 8'hfd ;
            rom[28161] = 8'hdc ;
            rom[28162] = 8'h10 ;
            rom[28163] = 8'he2 ;
            rom[28164] = 8'h1a ;
            rom[28165] = 8'h1e ;
            rom[28166] = 8'h2e ;
            rom[28167] = 8'h1c ;
            rom[28168] = 8'hd6 ;
            rom[28169] = 8'hc6 ;
            rom[28170] = 8'h0e ;
            rom[28171] = 8'hdf ;
            rom[28172] = 8'hef ;
            rom[28173] = 8'hfd ;
            rom[28174] = 8'h0f ;
            rom[28175] = 8'hfc ;
            rom[28176] = 8'he6 ;
            rom[28177] = 8'h09 ;
            rom[28178] = 8'hd5 ;
            rom[28179] = 8'hb1 ;
            rom[28180] = 8'hca ;
            rom[28181] = 8'h05 ;
            rom[28182] = 8'h1e ;
            rom[28183] = 8'hec ;
            rom[28184] = 8'hde ;
            rom[28185] = 8'hc2 ;
            rom[28186] = 8'hff ;
            rom[28187] = 8'h20 ;
            rom[28188] = 8'h34 ;
            rom[28189] = 8'hff ;
            rom[28190] = 8'hed ;
            rom[28191] = 8'hf8 ;
            rom[28192] = 8'hf4 ;
            rom[28193] = 8'h1d ;
            rom[28194] = 8'h0b ;
            rom[28195] = 8'hf4 ;
            rom[28196] = 8'hff ;
            rom[28197] = 8'hfe ;
            rom[28198] = 8'h27 ;
            rom[28199] = 8'hdf ;
            rom[28200] = 8'h13 ;
            rom[28201] = 8'h0b ;
            rom[28202] = 8'h07 ;
            rom[28203] = 8'he4 ;
            rom[28204] = 8'hff ;
            rom[28205] = 8'he8 ;
            rom[28206] = 8'h11 ;
            rom[28207] = 8'hfb ;
            rom[28208] = 8'h05 ;
            rom[28209] = 8'h0a ;
            rom[28210] = 8'h13 ;
            rom[28211] = 8'he7 ;
            rom[28212] = 8'hf8 ;
            rom[28213] = 8'hff ;
            rom[28214] = 8'h00 ;
            rom[28215] = 8'h0f ;
            rom[28216] = 8'he8 ;
            rom[28217] = 8'he0 ;
            rom[28218] = 8'h02 ;
            rom[28219] = 8'hdb ;
            rom[28220] = 8'h07 ;
            rom[28221] = 8'h1b ;
            rom[28222] = 8'h04 ;
            rom[28223] = 8'hfd ;
            rom[28224] = 8'h1a ;
            rom[28225] = 8'h13 ;
            rom[28226] = 8'hce ;
            rom[28227] = 8'hef ;
            rom[28228] = 8'hf4 ;
            rom[28229] = 8'he7 ;
            rom[28230] = 8'hf7 ;
            rom[28231] = 8'h07 ;
            rom[28232] = 8'h01 ;
            rom[28233] = 8'h1c ;
            rom[28234] = 8'h13 ;
            rom[28235] = 8'h23 ;
            rom[28236] = 8'he2 ;
            rom[28237] = 8'hf4 ;
            rom[28238] = 8'h0f ;
            rom[28239] = 8'h21 ;
            rom[28240] = 8'hf9 ;
            rom[28241] = 8'h10 ;
            rom[28242] = 8'h1e ;
            rom[28243] = 8'hea ;
            rom[28244] = 8'h08 ;
            rom[28245] = 8'h12 ;
            rom[28246] = 8'hf6 ;
            rom[28247] = 8'h1e ;
            rom[28248] = 8'h06 ;
            rom[28249] = 8'hfd ;
            rom[28250] = 8'h1a ;
            rom[28251] = 8'h1d ;
            rom[28252] = 8'hf3 ;
            rom[28253] = 8'hf4 ;
            rom[28254] = 8'h03 ;
            rom[28255] = 8'hfa ;
            rom[28256] = 8'hb3 ;
            rom[28257] = 8'hef ;
            rom[28258] = 8'hfc ;
            rom[28259] = 8'hf1 ;
            rom[28260] = 8'hf8 ;
            rom[28261] = 8'hd8 ;
            rom[28262] = 8'he5 ;
            rom[28263] = 8'h0a ;
            rom[28264] = 8'h19 ;
            rom[28265] = 8'h18 ;
            rom[28266] = 8'h17 ;
            rom[28267] = 8'h0d ;
            rom[28268] = 8'h04 ;
            rom[28269] = 8'h13 ;
            rom[28270] = 8'h0b ;
            rom[28271] = 8'h03 ;
            rom[28272] = 8'hfd ;
            rom[28273] = 8'h20 ;
            rom[28274] = 8'h1b ;
            rom[28275] = 8'h11 ;
            rom[28276] = 8'hf5 ;
            rom[28277] = 8'h05 ;
            rom[28278] = 8'h17 ;
            rom[28279] = 8'h1b ;
            rom[28280] = 8'h05 ;
            rom[28281] = 8'hc9 ;
            rom[28282] = 8'hfb ;
            rom[28283] = 8'h15 ;
            rom[28284] = 8'hf9 ;
            rom[28285] = 8'hfc ;
            rom[28286] = 8'h0a ;
            rom[28287] = 8'hc7 ;
            rom[28288] = 8'hf8 ;
            rom[28289] = 8'hff ;
            rom[28290] = 8'h04 ;
            rom[28291] = 8'he9 ;
            rom[28292] = 8'h09 ;
            rom[28293] = 8'hec ;
            rom[28294] = 8'h0b ;
            rom[28295] = 8'h15 ;
            rom[28296] = 8'h00 ;
            rom[28297] = 8'hd9 ;
            rom[28298] = 8'h04 ;
            rom[28299] = 8'hf6 ;
            rom[28300] = 8'hf9 ;
            rom[28301] = 8'hd7 ;
            rom[28302] = 8'hf0 ;
            rom[28303] = 8'h05 ;
            rom[28304] = 8'h0d ;
            rom[28305] = 8'he5 ;
            rom[28306] = 8'h07 ;
            rom[28307] = 8'h05 ;
            rom[28308] = 8'he8 ;
            rom[28309] = 8'hfb ;
            rom[28310] = 8'hfb ;
            rom[28311] = 8'h18 ;
            rom[28312] = 8'hf2 ;
            rom[28313] = 8'he8 ;
            rom[28314] = 8'h1e ;
            rom[28315] = 8'he1 ;
            rom[28316] = 8'h04 ;
            rom[28317] = 8'hfa ;
            rom[28318] = 8'hf7 ;
            rom[28319] = 8'h0b ;
            rom[28320] = 8'h0f ;
            rom[28321] = 8'h37 ;
            rom[28322] = 8'h0d ;
            rom[28323] = 8'hfd ;
            rom[28324] = 8'hf5 ;
            rom[28325] = 8'hfd ;
            rom[28326] = 8'hd5 ;
            rom[28327] = 8'h1a ;
            rom[28328] = 8'heb ;
            rom[28329] = 8'hf5 ;
            rom[28330] = 8'h09 ;
            rom[28331] = 8'h11 ;
            rom[28332] = 8'he0 ;
            rom[28333] = 8'h0f ;
            rom[28334] = 8'hfa ;
            rom[28335] = 8'hec ;
            rom[28336] = 8'h13 ;
            rom[28337] = 8'h06 ;
            rom[28338] = 8'hec ;
            rom[28339] = 8'h00 ;
            rom[28340] = 8'hfb ;
            rom[28341] = 8'h07 ;
            rom[28342] = 8'h18 ;
            rom[28343] = 8'hf5 ;
            rom[28344] = 8'hf9 ;
            rom[28345] = 8'hfa ;
            rom[28346] = 8'h11 ;
            rom[28347] = 8'h03 ;
            rom[28348] = 8'hf7 ;
            rom[28349] = 8'h09 ;
            rom[28350] = 8'h24 ;
            rom[28351] = 8'hb3 ;
            rom[28352] = 8'hd8 ;
            rom[28353] = 8'hef ;
            rom[28354] = 8'hf2 ;
            rom[28355] = 8'hfd ;
            rom[28356] = 8'hdb ;
            rom[28357] = 8'hf8 ;
            rom[28358] = 8'hd9 ;
            rom[28359] = 8'hfe ;
            rom[28360] = 8'h1a ;
            rom[28361] = 8'h0a ;
            rom[28362] = 8'h0d ;
            rom[28363] = 8'hea ;
            rom[28364] = 8'h03 ;
            rom[28365] = 8'h11 ;
            rom[28366] = 8'hf9 ;
            rom[28367] = 8'h00 ;
            rom[28368] = 8'hec ;
            rom[28369] = 8'hef ;
            rom[28370] = 8'h05 ;
            rom[28371] = 8'hff ;
            rom[28372] = 8'h06 ;
            rom[28373] = 8'he9 ;
            rom[28374] = 8'h15 ;
            rom[28375] = 8'he2 ;
            rom[28376] = 8'h03 ;
            rom[28377] = 8'h14 ;
            rom[28378] = 8'hee ;
            rom[28379] = 8'hfd ;
            rom[28380] = 8'hed ;
            rom[28381] = 8'hf9 ;
            rom[28382] = 8'hdf ;
            rom[28383] = 8'h1e ;
            rom[28384] = 8'h0d ;
            rom[28385] = 8'hef ;
            rom[28386] = 8'hf5 ;
            rom[28387] = 8'hf2 ;
            rom[28388] = 8'h08 ;
            rom[28389] = 8'h06 ;
            rom[28390] = 8'hf8 ;
            rom[28391] = 8'hc3 ;
            rom[28392] = 8'hdd ;
            rom[28393] = 8'hc5 ;
            rom[28394] = 8'hd8 ;
            rom[28395] = 8'hf4 ;
            rom[28396] = 8'hf5 ;
            rom[28397] = 8'hec ;
            rom[28398] = 8'h10 ;
            rom[28399] = 8'hda ;
            rom[28400] = 8'hf9 ;
            rom[28401] = 8'he2 ;
            rom[28402] = 8'hf1 ;
            rom[28403] = 8'hea ;
            rom[28404] = 8'hf9 ;
            rom[28405] = 8'he2 ;
            rom[28406] = 8'he0 ;
            rom[28407] = 8'he0 ;
            rom[28408] = 8'hf9 ;
            rom[28409] = 8'hd1 ;
            rom[28410] = 8'hf9 ;
            rom[28411] = 8'h16 ;
            rom[28412] = 8'he1 ;
            rom[28413] = 8'hd1 ;
            rom[28414] = 8'h23 ;
            rom[28415] = 8'h2c ;
            rom[28416] = 8'hee ;
            rom[28417] = 8'h0e ;
            rom[28418] = 8'hf7 ;
            rom[28419] = 8'h11 ;
            rom[28420] = 8'h05 ;
            rom[28421] = 8'h00 ;
            rom[28422] = 8'hdc ;
            rom[28423] = 8'h30 ;
            rom[28424] = 8'hec ;
            rom[28425] = 8'hf6 ;
            rom[28426] = 8'h14 ;
            rom[28427] = 8'he6 ;
            rom[28428] = 8'h00 ;
            rom[28429] = 8'hd2 ;
            rom[28430] = 8'h08 ;
            rom[28431] = 8'hdc ;
            rom[28432] = 8'hf3 ;
            rom[28433] = 8'hfc ;
            rom[28434] = 8'h0c ;
            rom[28435] = 8'h14 ;
            rom[28436] = 8'h01 ;
            rom[28437] = 8'hfe ;
            rom[28438] = 8'h02 ;
            rom[28439] = 8'h21 ;
            rom[28440] = 8'hf3 ;
            rom[28441] = 8'h18 ;
            rom[28442] = 8'h01 ;
            rom[28443] = 8'h0c ;
            rom[28444] = 8'hd8 ;
            rom[28445] = 8'h08 ;
            rom[28446] = 8'h2f ;
            rom[28447] = 8'h0a ;
            rom[28448] = 8'hc0 ;
            rom[28449] = 8'hf1 ;
            rom[28450] = 8'h0e ;
            rom[28451] = 8'h2a ;
            rom[28452] = 8'h08 ;
            rom[28453] = 8'h29 ;
            rom[28454] = 8'h04 ;
            rom[28455] = 8'h0b ;
            rom[28456] = 8'h08 ;
            rom[28457] = 8'hf0 ;
            rom[28458] = 8'hf7 ;
            rom[28459] = 8'h09 ;
            rom[28460] = 8'he7 ;
            rom[28461] = 8'hdf ;
            rom[28462] = 8'he7 ;
            rom[28463] = 8'h18 ;
            rom[28464] = 8'h1d ;
            rom[28465] = 8'h1a ;
            rom[28466] = 8'h0b ;
            rom[28467] = 8'hf0 ;
            rom[28468] = 8'hec ;
            rom[28469] = 8'h0e ;
            rom[28470] = 8'h1b ;
            rom[28471] = 8'hf3 ;
            rom[28472] = 8'h0e ;
            rom[28473] = 8'h0a ;
            rom[28474] = 8'hf9 ;
            rom[28475] = 8'h21 ;
            rom[28476] = 8'hf8 ;
            rom[28477] = 8'h06 ;
            rom[28478] = 8'hee ;
            rom[28479] = 8'hf7 ;
            rom[28480] = 8'hfb ;
            rom[28481] = 8'hef ;
            rom[28482] = 8'hbb ;
            rom[28483] = 8'h02 ;
            rom[28484] = 8'h1e ;
            rom[28485] = 8'h00 ;
            rom[28486] = 8'hf0 ;
            rom[28487] = 8'h00 ;
            rom[28488] = 8'hf7 ;
            rom[28489] = 8'h01 ;
            rom[28490] = 8'hed ;
            rom[28491] = 8'h25 ;
            rom[28492] = 8'hfc ;
            rom[28493] = 8'hf9 ;
            rom[28494] = 8'hd6 ;
            rom[28495] = 8'hd3 ;
            rom[28496] = 8'hff ;
            rom[28497] = 8'hfa ;
            rom[28498] = 8'h0e ;
            rom[28499] = 8'h02 ;
            rom[28500] = 8'hf4 ;
            rom[28501] = 8'h20 ;
            rom[28502] = 8'h08 ;
            rom[28503] = 8'hee ;
            rom[28504] = 8'h15 ;
            rom[28505] = 8'h21 ;
            rom[28506] = 8'h1e ;
            rom[28507] = 8'he8 ;
            rom[28508] = 8'h0c ;
            rom[28509] = 8'hf9 ;
            rom[28510] = 8'h09 ;
            rom[28511] = 8'hf6 ;
            rom[28512] = 8'hf2 ;
            rom[28513] = 8'h11 ;
            rom[28514] = 8'hdf ;
            rom[28515] = 8'he5 ;
            rom[28516] = 8'hd8 ;
            rom[28517] = 8'hf3 ;
            rom[28518] = 8'hfd ;
            rom[28519] = 8'hf6 ;
            rom[28520] = 8'hf3 ;
            rom[28521] = 8'he0 ;
            rom[28522] = 8'hce ;
            rom[28523] = 8'h03 ;
            rom[28524] = 8'hee ;
            rom[28525] = 8'hee ;
            rom[28526] = 8'h0b ;
            rom[28527] = 8'hdb ;
            rom[28528] = 8'h02 ;
            rom[28529] = 8'hfa ;
            rom[28530] = 8'h14 ;
            rom[28531] = 8'he1 ;
            rom[28532] = 8'hf9 ;
            rom[28533] = 8'hc7 ;
            rom[28534] = 8'h0b ;
            rom[28535] = 8'hec ;
            rom[28536] = 8'he2 ;
            rom[28537] = 8'h04 ;
            rom[28538] = 8'hec ;
            rom[28539] = 8'h26 ;
            rom[28540] = 8'hf2 ;
            rom[28541] = 8'hc6 ;
            rom[28542] = 8'h1e ;
            rom[28543] = 8'h0b ;
            rom[28544] = 8'h06 ;
            rom[28545] = 8'hf3 ;
            rom[28546] = 8'he7 ;
            rom[28547] = 8'he1 ;
            rom[28548] = 8'hf4 ;
            rom[28549] = 8'hfc ;
            rom[28550] = 8'hef ;
            rom[28551] = 8'h02 ;
            rom[28552] = 8'h30 ;
            rom[28553] = 8'hda ;
            rom[28554] = 8'h02 ;
            rom[28555] = 8'hf0 ;
            rom[28556] = 8'hd4 ;
            rom[28557] = 8'h19 ;
            rom[28558] = 8'h24 ;
            rom[28559] = 8'he0 ;
            rom[28560] = 8'hf8 ;
            rom[28561] = 8'hef ;
            rom[28562] = 8'hf7 ;
            rom[28563] = 8'hf9 ;
            rom[28564] = 8'hd5 ;
            rom[28565] = 8'hf3 ;
            rom[28566] = 8'hf6 ;
            rom[28567] = 8'hf7 ;
            rom[28568] = 8'hfb ;
            rom[28569] = 8'h13 ;
            rom[28570] = 8'h07 ;
            rom[28571] = 8'h20 ;
            rom[28572] = 8'h16 ;
            rom[28573] = 8'h0c ;
            rom[28574] = 8'hc7 ;
            rom[28575] = 8'hdf ;
            rom[28576] = 8'h02 ;
            rom[28577] = 8'hed ;
            rom[28578] = 8'h0a ;
            rom[28579] = 8'hef ;
            rom[28580] = 8'he6 ;
            rom[28581] = 8'he9 ;
            rom[28582] = 8'h00 ;
            rom[28583] = 8'hf5 ;
            rom[28584] = 8'hfd ;
            rom[28585] = 8'hf1 ;
            rom[28586] = 8'h0b ;
            rom[28587] = 8'hf6 ;
            rom[28588] = 8'hf6 ;
            rom[28589] = 8'hf2 ;
            rom[28590] = 8'hf2 ;
            rom[28591] = 8'hf6 ;
            rom[28592] = 8'h0d ;
            rom[28593] = 8'h04 ;
            rom[28594] = 8'hf7 ;
            rom[28595] = 8'h18 ;
            rom[28596] = 8'he4 ;
            rom[28597] = 8'hea ;
            rom[28598] = 8'hdf ;
            rom[28599] = 8'h18 ;
            rom[28600] = 8'h02 ;
            rom[28601] = 8'hfd ;
            rom[28602] = 8'he2 ;
            rom[28603] = 8'hb5 ;
            rom[28604] = 8'he9 ;
            rom[28605] = 8'h0c ;
            rom[28606] = 8'hf5 ;
            rom[28607] = 8'hcd ;
            rom[28608] = 8'h0a ;
            rom[28609] = 8'h18 ;
            rom[28610] = 8'h0e ;
            rom[28611] = 8'hed ;
            rom[28612] = 8'hf6 ;
            rom[28613] = 8'h16 ;
            rom[28614] = 8'h04 ;
            rom[28615] = 8'hf4 ;
            rom[28616] = 8'he7 ;
            rom[28617] = 8'hee ;
            rom[28618] = 8'h08 ;
            rom[28619] = 8'hc9 ;
            rom[28620] = 8'hf7 ;
            rom[28621] = 8'hfb ;
            rom[28622] = 8'h0b ;
            rom[28623] = 8'hd6 ;
            rom[28624] = 8'h14 ;
            rom[28625] = 8'hfd ;
            rom[28626] = 8'h0c ;
            rom[28627] = 8'hf0 ;
            rom[28628] = 8'h00 ;
            rom[28629] = 8'hf0 ;
            rom[28630] = 8'hf3 ;
            rom[28631] = 8'h2c ;
            rom[28632] = 8'hee ;
            rom[28633] = 8'hf7 ;
            rom[28634] = 8'hf3 ;
            rom[28635] = 8'hfb ;
            rom[28636] = 8'h12 ;
            rom[28637] = 8'hf3 ;
            rom[28638] = 8'hc8 ;
            rom[28639] = 8'hf4 ;
            rom[28640] = 8'hf3 ;
            rom[28641] = 8'hee ;
            rom[28642] = 8'hcc ;
            rom[28643] = 8'hf5 ;
            rom[28644] = 8'he4 ;
            rom[28645] = 8'he0 ;
            rom[28646] = 8'hf4 ;
            rom[28647] = 8'he6 ;
            rom[28648] = 8'h03 ;
            rom[28649] = 8'hfc ;
            rom[28650] = 8'hfd ;
            rom[28651] = 8'hfe ;
            rom[28652] = 8'h11 ;
            rom[28653] = 8'hcb ;
            rom[28654] = 8'he1 ;
            rom[28655] = 8'hf1 ;
            rom[28656] = 8'hde ;
            rom[28657] = 8'hfb ;
            rom[28658] = 8'h06 ;
            rom[28659] = 8'h1b ;
            rom[28660] = 8'hd4 ;
            rom[28661] = 8'h0a ;
            rom[28662] = 8'hfe ;
            rom[28663] = 8'hef ;
            rom[28664] = 8'hf7 ;
            rom[28665] = 8'hf8 ;
            rom[28666] = 8'hea ;
            rom[28667] = 8'he3 ;
            rom[28668] = 8'hef ;
            rom[28669] = 8'h0d ;
            rom[28670] = 8'h03 ;
            rom[28671] = 8'he2 ;
            rom[28672] = 8'hf1 ;
            rom[28673] = 8'h0c ;
            rom[28674] = 8'hda ;
            rom[28675] = 8'h26 ;
            rom[28676] = 8'h37 ;
            rom[28677] = 8'hef ;
            rom[28678] = 8'hcf ;
            rom[28679] = 8'h0f ;
            rom[28680] = 8'he9 ;
            rom[28681] = 8'h01 ;
            rom[28682] = 8'h1a ;
            rom[28683] = 8'hbc ;
            rom[28684] = 8'hce ;
            rom[28685] = 8'hd8 ;
            rom[28686] = 8'h0f ;
            rom[28687] = 8'he6 ;
            rom[28688] = 8'hdc ;
            rom[28689] = 8'hff ;
            rom[28690] = 8'h08 ;
            rom[28691] = 8'hf8 ;
            rom[28692] = 8'h0d ;
            rom[28693] = 8'he3 ;
            rom[28694] = 8'h0e ;
            rom[28695] = 8'h05 ;
            rom[28696] = 8'hf8 ;
            rom[28697] = 8'hde ;
            rom[28698] = 8'h16 ;
            rom[28699] = 8'hf6 ;
            rom[28700] = 8'h11 ;
            rom[28701] = 8'he4 ;
            rom[28702] = 8'hf8 ;
            rom[28703] = 8'hff ;
            rom[28704] = 8'hfb ;
            rom[28705] = 8'hff ;
            rom[28706] = 8'hf3 ;
            rom[28707] = 8'h15 ;
            rom[28708] = 8'hd5 ;
            rom[28709] = 8'hd7 ;
            rom[28710] = 8'hb1 ;
            rom[28711] = 8'h0d ;
            rom[28712] = 8'he1 ;
            rom[28713] = 8'hf6 ;
            rom[28714] = 8'h00 ;
            rom[28715] = 8'h1b ;
            rom[28716] = 8'he4 ;
            rom[28717] = 8'hc9 ;
            rom[28718] = 8'he4 ;
            rom[28719] = 8'h1b ;
            rom[28720] = 8'h23 ;
            rom[28721] = 8'hf2 ;
            rom[28722] = 8'h03 ;
            rom[28723] = 8'hf5 ;
            rom[28724] = 8'hb1 ;
            rom[28725] = 8'h16 ;
            rom[28726] = 8'h09 ;
            rom[28727] = 8'hf9 ;
            rom[28728] = 8'hff ;
            rom[28729] = 8'hf1 ;
            rom[28730] = 8'h18 ;
            rom[28731] = 8'h00 ;
            rom[28732] = 8'hfb ;
            rom[28733] = 8'hfa ;
            rom[28734] = 8'h0c ;
            rom[28735] = 8'hed ;
            rom[28736] = 8'hf2 ;
            rom[28737] = 8'h09 ;
            rom[28738] = 8'hde ;
            rom[28739] = 8'h12 ;
            rom[28740] = 8'hfd ;
            rom[28741] = 8'hff ;
            rom[28742] = 8'hdd ;
            rom[28743] = 8'hf6 ;
            rom[28744] = 8'hf2 ;
            rom[28745] = 8'hf4 ;
            rom[28746] = 8'hf8 ;
            rom[28747] = 8'hec ;
            rom[28748] = 8'he2 ;
            rom[28749] = 8'hc9 ;
            rom[28750] = 8'hd2 ;
            rom[28751] = 8'hed ;
            rom[28752] = 8'h05 ;
            rom[28753] = 8'he2 ;
            rom[28754] = 8'h13 ;
            rom[28755] = 8'hd5 ;
            rom[28756] = 8'h0e ;
            rom[28757] = 8'h0c ;
            rom[28758] = 8'hd0 ;
            rom[28759] = 8'h0b ;
            rom[28760] = 8'h04 ;
            rom[28761] = 8'h1e ;
            rom[28762] = 8'h0b ;
            rom[28763] = 8'h1a ;
            rom[28764] = 8'hfa ;
            rom[28765] = 8'hf2 ;
            rom[28766] = 8'hea ;
            rom[28767] = 8'he5 ;
            rom[28768] = 8'hd1 ;
            rom[28769] = 8'hfc ;
            rom[28770] = 8'hfd ;
            rom[28771] = 8'he2 ;
            rom[28772] = 8'heb ;
            rom[28773] = 8'hfa ;
            rom[28774] = 8'hf9 ;
            rom[28775] = 8'he1 ;
            rom[28776] = 8'hed ;
            rom[28777] = 8'h0a ;
            rom[28778] = 8'h02 ;
            rom[28779] = 8'he3 ;
            rom[28780] = 8'h1b ;
            rom[28781] = 8'hfc ;
            rom[28782] = 8'hf0 ;
            rom[28783] = 8'h1a ;
            rom[28784] = 8'he6 ;
            rom[28785] = 8'hee ;
            rom[28786] = 8'h08 ;
            rom[28787] = 8'hff ;
            rom[28788] = 8'he2 ;
            rom[28789] = 8'he2 ;
            rom[28790] = 8'hf0 ;
            rom[28791] = 8'h05 ;
            rom[28792] = 8'h00 ;
            rom[28793] = 8'he2 ;
            rom[28794] = 8'hf2 ;
            rom[28795] = 8'h04 ;
            rom[28796] = 8'hf0 ;
            rom[28797] = 8'h20 ;
            rom[28798] = 8'h04 ;
            rom[28799] = 8'h01 ;
            rom[28800] = 8'h0c ;
            rom[28801] = 8'ha8 ;
            rom[28802] = 8'h0f ;
            rom[28803] = 8'hdd ;
            rom[28804] = 8'hfb ;
            rom[28805] = 8'h18 ;
            rom[28806] = 8'hc5 ;
            rom[28807] = 8'hfb ;
            rom[28808] = 8'hde ;
            rom[28809] = 8'hf7 ;
            rom[28810] = 8'h1e ;
            rom[28811] = 8'hf1 ;
            rom[28812] = 8'h05 ;
            rom[28813] = 8'h07 ;
            rom[28814] = 8'h24 ;
            rom[28815] = 8'h1e ;
            rom[28816] = 8'hf0 ;
            rom[28817] = 8'hfb ;
            rom[28818] = 8'hcc ;
            rom[28819] = 8'hdf ;
            rom[28820] = 8'he8 ;
            rom[28821] = 8'hdf ;
            rom[28822] = 8'hfe ;
            rom[28823] = 8'hfc ;
            rom[28824] = 8'h03 ;
            rom[28825] = 8'hde ;
            rom[28826] = 8'hf2 ;
            rom[28827] = 8'h04 ;
            rom[28828] = 8'h1a ;
            rom[28829] = 8'hfe ;
            rom[28830] = 8'hda ;
            rom[28831] = 8'hfa ;
            rom[28832] = 8'h21 ;
            rom[28833] = 8'hf5 ;
            rom[28834] = 8'hd9 ;
            rom[28835] = 8'hea ;
            rom[28836] = 8'hff ;
            rom[28837] = 8'hee ;
            rom[28838] = 8'h17 ;
            rom[28839] = 8'hd8 ;
            rom[28840] = 8'h06 ;
            rom[28841] = 8'hdf ;
            rom[28842] = 8'h04 ;
            rom[28843] = 8'hf2 ;
            rom[28844] = 8'hfb ;
            rom[28845] = 8'hda ;
            rom[28846] = 8'hf3 ;
            rom[28847] = 8'hed ;
            rom[28848] = 8'h10 ;
            rom[28849] = 8'hff ;
            rom[28850] = 8'hdf ;
            rom[28851] = 8'h03 ;
            rom[28852] = 8'h13 ;
            rom[28853] = 8'hd8 ;
            rom[28854] = 8'h21 ;
            rom[28855] = 8'he5 ;
            rom[28856] = 8'h1c ;
            rom[28857] = 8'h15 ;
            rom[28858] = 8'hf2 ;
            rom[28859] = 8'hfe ;
            rom[28860] = 8'h12 ;
            rom[28861] = 8'h1a ;
            rom[28862] = 8'hee ;
            rom[28863] = 8'h02 ;
            rom[28864] = 8'he8 ;
            rom[28865] = 8'h00 ;
            rom[28866] = 8'h1d ;
            rom[28867] = 8'hff ;
            rom[28868] = 8'hc0 ;
            rom[28869] = 8'h00 ;
            rom[28870] = 8'he8 ;
            rom[28871] = 8'h13 ;
            rom[28872] = 8'hf5 ;
            rom[28873] = 8'h21 ;
            rom[28874] = 8'h14 ;
            rom[28875] = 8'hfe ;
            rom[28876] = 8'hfe ;
            rom[28877] = 8'hf7 ;
            rom[28878] = 8'h08 ;
            rom[28879] = 8'h1a ;
            rom[28880] = 8'h08 ;
            rom[28881] = 8'h16 ;
            rom[28882] = 8'hcc ;
            rom[28883] = 8'hee ;
            rom[28884] = 8'hfa ;
            rom[28885] = 8'he5 ;
            rom[28886] = 8'hd5 ;
            rom[28887] = 8'h1a ;
            rom[28888] = 8'he2 ;
            rom[28889] = 8'hf6 ;
            rom[28890] = 8'he2 ;
            rom[28891] = 8'h03 ;
            rom[28892] = 8'h29 ;
            rom[28893] = 8'he7 ;
            rom[28894] = 8'h16 ;
            rom[28895] = 8'hf9 ;
            rom[28896] = 8'hed ;
            rom[28897] = 8'h0a ;
            rom[28898] = 8'hfb ;
            rom[28899] = 8'hf4 ;
            rom[28900] = 8'hd7 ;
            rom[28901] = 8'hee ;
            rom[28902] = 8'h01 ;
            rom[28903] = 8'h1f ;
            rom[28904] = 8'hff ;
            rom[28905] = 8'h09 ;
            rom[28906] = 8'hd7 ;
            rom[28907] = 8'hfd ;
            rom[28908] = 8'hf6 ;
            rom[28909] = 8'h09 ;
            rom[28910] = 8'h20 ;
            rom[28911] = 8'h1e ;
            rom[28912] = 8'h17 ;
            rom[28913] = 8'h08 ;
            rom[28914] = 8'hfb ;
            rom[28915] = 8'h19 ;
            rom[28916] = 8'h08 ;
            rom[28917] = 8'h17 ;
            rom[28918] = 8'he3 ;
            rom[28919] = 8'h1d ;
            rom[28920] = 8'hf9 ;
            rom[28921] = 8'h01 ;
            rom[28922] = 8'hf6 ;
            rom[28923] = 8'h08 ;
            rom[28924] = 8'hf2 ;
            rom[28925] = 8'h12 ;
            rom[28926] = 8'hd6 ;
            rom[28927] = 8'hf2 ;
            rom[28928] = 8'h16 ;
            rom[28929] = 8'h21 ;
            rom[28930] = 8'h00 ;
            rom[28931] = 8'hf6 ;
            rom[28932] = 8'h08 ;
            rom[28933] = 8'h00 ;
            rom[28934] = 8'hfc ;
            rom[28935] = 8'h1a ;
            rom[28936] = 8'h01 ;
            rom[28937] = 8'hd7 ;
            rom[28938] = 8'h10 ;
            rom[28939] = 8'he8 ;
            rom[28940] = 8'hf2 ;
            rom[28941] = 8'hfd ;
            rom[28942] = 8'h04 ;
            rom[28943] = 8'hfd ;
            rom[28944] = 8'h06 ;
            rom[28945] = 8'he3 ;
            rom[28946] = 8'h02 ;
            rom[28947] = 8'h09 ;
            rom[28948] = 8'h05 ;
            rom[28949] = 8'h1f ;
            rom[28950] = 8'hdd ;
            rom[28951] = 8'h1d ;
            rom[28952] = 8'he6 ;
            rom[28953] = 8'hbd ;
            rom[28954] = 8'h0b ;
            rom[28955] = 8'hd2 ;
            rom[28956] = 8'h04 ;
            rom[28957] = 8'h0b ;
            rom[28958] = 8'hf1 ;
            rom[28959] = 8'hf9 ;
            rom[28960] = 8'h00 ;
            rom[28961] = 8'h12 ;
            rom[28962] = 8'hfb ;
            rom[28963] = 8'h0d ;
            rom[28964] = 8'he5 ;
            rom[28965] = 8'h10 ;
            rom[28966] = 8'hec ;
            rom[28967] = 8'h08 ;
            rom[28968] = 8'h0b ;
            rom[28969] = 8'h05 ;
            rom[28970] = 8'h11 ;
            rom[28971] = 8'h12 ;
            rom[28972] = 8'h02 ;
            rom[28973] = 8'hfe ;
            rom[28974] = 8'h08 ;
            rom[28975] = 8'hf3 ;
            rom[28976] = 8'h20 ;
            rom[28977] = 8'h0f ;
            rom[28978] = 8'hef ;
            rom[28979] = 8'hc3 ;
            rom[28980] = 8'hef ;
            rom[28981] = 8'hec ;
            rom[28982] = 8'h18 ;
            rom[28983] = 8'h0b ;
            rom[28984] = 8'h2a ;
            rom[28985] = 8'ha9 ;
            rom[28986] = 8'h02 ;
            rom[28987] = 8'h13 ;
            rom[28988] = 8'h29 ;
            rom[28989] = 8'he6 ;
            rom[28990] = 8'h0b ;
            rom[28991] = 8'hbf ;
            rom[28992] = 8'h12 ;
            rom[28993] = 8'h04 ;
            rom[28994] = 8'he3 ;
            rom[28995] = 8'h05 ;
            rom[28996] = 8'hd5 ;
            rom[28997] = 8'h1a ;
            rom[28998] = 8'hdf ;
            rom[28999] = 8'hf1 ;
            rom[29000] = 8'h22 ;
            rom[29001] = 8'h04 ;
            rom[29002] = 8'hef ;
            rom[29003] = 8'h14 ;
            rom[29004] = 8'hb5 ;
            rom[29005] = 8'h09 ;
            rom[29006] = 8'he9 ;
            rom[29007] = 8'hfc ;
            rom[29008] = 8'h0b ;
            rom[29009] = 8'h03 ;
            rom[29010] = 8'hfe ;
            rom[29011] = 8'he4 ;
            rom[29012] = 8'h2b ;
            rom[29013] = 8'hfe ;
            rom[29014] = 8'hd4 ;
            rom[29015] = 8'hee ;
            rom[29016] = 8'h0a ;
            rom[29017] = 8'h1e ;
            rom[29018] = 8'h04 ;
            rom[29019] = 8'hf2 ;
            rom[29020] = 8'h09 ;
            rom[29021] = 8'h08 ;
            rom[29022] = 8'hff ;
            rom[29023] = 8'h14 ;
            rom[29024] = 8'hd7 ;
            rom[29025] = 8'h23 ;
            rom[29026] = 8'hf7 ;
            rom[29027] = 8'h04 ;
            rom[29028] = 8'hef ;
            rom[29029] = 8'hf0 ;
            rom[29030] = 8'h22 ;
            rom[29031] = 8'he0 ;
            rom[29032] = 8'he0 ;
            rom[29033] = 8'h0b ;
            rom[29034] = 8'he9 ;
            rom[29035] = 8'hf4 ;
            rom[29036] = 8'h17 ;
            rom[29037] = 8'h18 ;
            rom[29038] = 8'h05 ;
            rom[29039] = 8'hf0 ;
            rom[29040] = 8'hdf ;
            rom[29041] = 8'h06 ;
            rom[29042] = 8'hec ;
            rom[29043] = 8'h13 ;
            rom[29044] = 8'h1d ;
            rom[29045] = 8'h0d ;
            rom[29046] = 8'hff ;
            rom[29047] = 8'h09 ;
            rom[29048] = 8'h03 ;
            rom[29049] = 8'h1d ;
            rom[29050] = 8'hd5 ;
            rom[29051] = 8'h06 ;
            rom[29052] = 8'h06 ;
            rom[29053] = 8'h12 ;
            rom[29054] = 8'h1b ;
            rom[29055] = 8'hf1 ;
            rom[29056] = 8'h13 ;
            rom[29057] = 8'he5 ;
            rom[29058] = 8'hde ;
            rom[29059] = 8'hf8 ;
            rom[29060] = 8'hfe ;
            rom[29061] = 8'h10 ;
            rom[29062] = 8'hf0 ;
            rom[29063] = 8'h03 ;
            rom[29064] = 8'h09 ;
            rom[29065] = 8'hec ;
            rom[29066] = 8'he9 ;
            rom[29067] = 8'h0f ;
            rom[29068] = 8'hde ;
            rom[29069] = 8'h23 ;
            rom[29070] = 8'h03 ;
            rom[29071] = 8'hf9 ;
            rom[29072] = 8'hfa ;
            rom[29073] = 8'hf9 ;
            rom[29074] = 8'hfd ;
            rom[29075] = 8'he5 ;
            rom[29076] = 8'hee ;
            rom[29077] = 8'hfc ;
            rom[29078] = 8'hff ;
            rom[29079] = 8'h13 ;
            rom[29080] = 8'hf5 ;
            rom[29081] = 8'hbf ;
            rom[29082] = 8'hf4 ;
            rom[29083] = 8'hed ;
            rom[29084] = 8'h02 ;
            rom[29085] = 8'h09 ;
            rom[29086] = 8'hb7 ;
            rom[29087] = 8'hff ;
            rom[29088] = 8'hf9 ;
            rom[29089] = 8'h22 ;
            rom[29090] = 8'hc5 ;
            rom[29091] = 8'h06 ;
            rom[29092] = 8'he7 ;
            rom[29093] = 8'h07 ;
            rom[29094] = 8'hf1 ;
            rom[29095] = 8'hcf ;
            rom[29096] = 8'hf6 ;
            rom[29097] = 8'hf7 ;
            rom[29098] = 8'h12 ;
            rom[29099] = 8'h12 ;
            rom[29100] = 8'h0c ;
            rom[29101] = 8'h11 ;
            rom[29102] = 8'he9 ;
            rom[29103] = 8'h12 ;
            rom[29104] = 8'hf3 ;
            rom[29105] = 8'heb ;
            rom[29106] = 8'hea ;
            rom[29107] = 8'hf0 ;
            rom[29108] = 8'h13 ;
            rom[29109] = 8'hea ;
            rom[29110] = 8'hf1 ;
            rom[29111] = 8'h0d ;
            rom[29112] = 8'h1e ;
            rom[29113] = 8'h12 ;
            rom[29114] = 8'hd7 ;
            rom[29115] = 8'hdd ;
            rom[29116] = 8'h16 ;
            rom[29117] = 8'h0a ;
            rom[29118] = 8'h12 ;
            rom[29119] = 8'hfd ;
            rom[29120] = 8'h03 ;
            rom[29121] = 8'h08 ;
            rom[29122] = 8'h06 ;
            rom[29123] = 8'hfc ;
            rom[29124] = 8'h02 ;
            rom[29125] = 8'h06 ;
            rom[29126] = 8'hce ;
            rom[29127] = 8'h02 ;
            rom[29128] = 8'he9 ;
            rom[29129] = 8'h11 ;
            rom[29130] = 8'h03 ;
            rom[29131] = 8'hf5 ;
            rom[29132] = 8'hd6 ;
            rom[29133] = 8'h0a ;
            rom[29134] = 8'h02 ;
            rom[29135] = 8'h23 ;
            rom[29136] = 8'h00 ;
            rom[29137] = 8'h13 ;
            rom[29138] = 8'he5 ;
            rom[29139] = 8'hec ;
            rom[29140] = 8'hee ;
            rom[29141] = 8'hf0 ;
            rom[29142] = 8'he3 ;
            rom[29143] = 8'h11 ;
            rom[29144] = 8'hd6 ;
            rom[29145] = 8'h1d ;
            rom[29146] = 8'hf9 ;
            rom[29147] = 8'hfb ;
            rom[29148] = 8'hd9 ;
            rom[29149] = 8'h1a ;
            rom[29150] = 8'h10 ;
            rom[29151] = 8'hf0 ;
            rom[29152] = 8'hc7 ;
            rom[29153] = 8'h1e ;
            rom[29154] = 8'hf1 ;
            rom[29155] = 8'h0e ;
            rom[29156] = 8'he3 ;
            rom[29157] = 8'hdc ;
            rom[29158] = 8'h01 ;
            rom[29159] = 8'h14 ;
            rom[29160] = 8'h19 ;
            rom[29161] = 8'h25 ;
            rom[29162] = 8'hf6 ;
            rom[29163] = 8'hfc ;
            rom[29164] = 8'h08 ;
            rom[29165] = 8'h02 ;
            rom[29166] = 8'hf0 ;
            rom[29167] = 8'h0d ;
            rom[29168] = 8'hfe ;
            rom[29169] = 8'h2c ;
            rom[29170] = 8'hf1 ;
            rom[29171] = 8'h11 ;
            rom[29172] = 8'h0c ;
            rom[29173] = 8'hf9 ;
            rom[29174] = 8'h0d ;
            rom[29175] = 8'hed ;
            rom[29176] = 8'hf9 ;
            rom[29177] = 8'h00 ;
            rom[29178] = 8'he7 ;
            rom[29179] = 8'he4 ;
            rom[29180] = 8'h07 ;
            rom[29181] = 8'h0d ;
            rom[29182] = 8'hcf ;
            rom[29183] = 8'hf8 ;
            rom[29184] = 8'h0e ;
            rom[29185] = 8'hfe ;
            rom[29186] = 8'hfd ;
            rom[29187] = 8'h0d ;
            rom[29188] = 8'hf8 ;
            rom[29189] = 8'hfe ;
            rom[29190] = 8'hed ;
            rom[29191] = 8'he0 ;
            rom[29192] = 8'h18 ;
            rom[29193] = 8'hf4 ;
            rom[29194] = 8'h0a ;
            rom[29195] = 8'h02 ;
            rom[29196] = 8'h09 ;
            rom[29197] = 8'h10 ;
            rom[29198] = 8'h11 ;
            rom[29199] = 8'h13 ;
            rom[29200] = 8'hc0 ;
            rom[29201] = 8'he3 ;
            rom[29202] = 8'h06 ;
            rom[29203] = 8'h00 ;
            rom[29204] = 8'hfe ;
            rom[29205] = 8'hd9 ;
            rom[29206] = 8'hf2 ;
            rom[29207] = 8'hf6 ;
            rom[29208] = 8'hfa ;
            rom[29209] = 8'h0e ;
            rom[29210] = 8'hd0 ;
            rom[29211] = 8'hb9 ;
            rom[29212] = 8'hf8 ;
            rom[29213] = 8'h00 ;
            rom[29214] = 8'hf5 ;
            rom[29215] = 8'hf7 ;
            rom[29216] = 8'hc3 ;
            rom[29217] = 8'heb ;
            rom[29218] = 8'hfb ;
            rom[29219] = 8'h00 ;
            rom[29220] = 8'he0 ;
            rom[29221] = 8'he3 ;
            rom[29222] = 8'h10 ;
            rom[29223] = 8'hd9 ;
            rom[29224] = 8'h0c ;
            rom[29225] = 8'he9 ;
            rom[29226] = 8'hfb ;
            rom[29227] = 8'hba ;
            rom[29228] = 8'h0b ;
            rom[29229] = 8'h10 ;
            rom[29230] = 8'hd8 ;
            rom[29231] = 8'hfd ;
            rom[29232] = 8'hf5 ;
            rom[29233] = 8'hff ;
            rom[29234] = 8'hf0 ;
            rom[29235] = 8'hfe ;
            rom[29236] = 8'hf2 ;
            rom[29237] = 8'hda ;
            rom[29238] = 8'he3 ;
            rom[29239] = 8'hf8 ;
            rom[29240] = 8'h01 ;
            rom[29241] = 8'hfa ;
            rom[29242] = 8'he2 ;
            rom[29243] = 8'hff ;
            rom[29244] = 8'he7 ;
            rom[29245] = 8'h11 ;
            rom[29246] = 8'hcc ;
            rom[29247] = 8'hec ;
            rom[29248] = 8'hfb ;
            rom[29249] = 8'he5 ;
            rom[29250] = 8'hf6 ;
            rom[29251] = 8'hfd ;
            rom[29252] = 8'hf6 ;
            rom[29253] = 8'h0a ;
            rom[29254] = 8'hf4 ;
            rom[29255] = 8'hc8 ;
            rom[29256] = 8'he8 ;
            rom[29257] = 8'h00 ;
            rom[29258] = 8'h1b ;
            rom[29259] = 8'h06 ;
            rom[29260] = 8'he1 ;
            rom[29261] = 8'hf9 ;
            rom[29262] = 8'hfa ;
            rom[29263] = 8'hce ;
            rom[29264] = 8'h18 ;
            rom[29265] = 8'h10 ;
            rom[29266] = 8'he6 ;
            rom[29267] = 8'h18 ;
            rom[29268] = 8'hf5 ;
            rom[29269] = 8'hdc ;
            rom[29270] = 8'hf4 ;
            rom[29271] = 8'hdb ;
            rom[29272] = 8'he8 ;
            rom[29273] = 8'hca ;
            rom[29274] = 8'hf8 ;
            rom[29275] = 8'hde ;
            rom[29276] = 8'hfa ;
            rom[29277] = 8'he9 ;
            rom[29278] = 8'h08 ;
            rom[29279] = 8'hf6 ;
            rom[29280] = 8'hf0 ;
            rom[29281] = 8'hf1 ;
            rom[29282] = 8'hee ;
            rom[29283] = 8'h0c ;
            rom[29284] = 8'hfc ;
            rom[29285] = 8'hf6 ;
            rom[29286] = 8'hf1 ;
            rom[29287] = 8'hdb ;
            rom[29288] = 8'h04 ;
            rom[29289] = 8'hec ;
            rom[29290] = 8'hfe ;
            rom[29291] = 8'h1d ;
            rom[29292] = 8'hdf ;
            rom[29293] = 8'hee ;
            rom[29294] = 8'hdc ;
            rom[29295] = 8'hf4 ;
            rom[29296] = 8'hef ;
            rom[29297] = 8'hea ;
            rom[29298] = 8'hfe ;
            rom[29299] = 8'hdf ;
            rom[29300] = 8'hc0 ;
            rom[29301] = 8'hf3 ;
            rom[29302] = 8'heb ;
            rom[29303] = 8'he0 ;
            rom[29304] = 8'h1c ;
            rom[29305] = 8'hf5 ;
            rom[29306] = 8'hfc ;
            rom[29307] = 8'hf0 ;
            rom[29308] = 8'hf2 ;
            rom[29309] = 8'hd2 ;
            rom[29310] = 8'hca ;
            rom[29311] = 8'hdf ;
            rom[29312] = 8'he0 ;
            rom[29313] = 8'hfb ;
            rom[29314] = 8'hf3 ;
            rom[29315] = 8'h07 ;
            rom[29316] = 8'hd8 ;
            rom[29317] = 8'h11 ;
            rom[29318] = 8'h15 ;
            rom[29319] = 8'h08 ;
            rom[29320] = 8'hf8 ;
            rom[29321] = 8'h2f ;
            rom[29322] = 8'hfe ;
            rom[29323] = 8'hfc ;
            rom[29324] = 8'h17 ;
            rom[29325] = 8'hf6 ;
            rom[29326] = 8'hf9 ;
            rom[29327] = 8'he2 ;
            rom[29328] = 8'h05 ;
            rom[29329] = 8'he0 ;
            rom[29330] = 8'hf9 ;
            rom[29331] = 8'h02 ;
            rom[29332] = 8'h10 ;
            rom[29333] = 8'hee ;
            rom[29334] = 8'hfb ;
            rom[29335] = 8'hf6 ;
            rom[29336] = 8'h0a ;
            rom[29337] = 8'h01 ;
            rom[29338] = 8'h09 ;
            rom[29339] = 8'hf3 ;
            rom[29340] = 8'he2 ;
            rom[29341] = 8'he8 ;
            rom[29342] = 8'hee ;
            rom[29343] = 8'hed ;
            rom[29344] = 8'hf0 ;
            rom[29345] = 8'h14 ;
            rom[29346] = 8'h0b ;
            rom[29347] = 8'hde ;
            rom[29348] = 8'h0b ;
            rom[29349] = 8'h20 ;
            rom[29350] = 8'h13 ;
            rom[29351] = 8'hfc ;
            rom[29352] = 8'he7 ;
            rom[29353] = 8'he3 ;
            rom[29354] = 8'h1c ;
            rom[29355] = 8'hfa ;
            rom[29356] = 8'heb ;
            rom[29357] = 8'hea ;
            rom[29358] = 8'h0e ;
            rom[29359] = 8'hea ;
            rom[29360] = 8'h00 ;
            rom[29361] = 8'hf1 ;
            rom[29362] = 8'h09 ;
            rom[29363] = 8'hea ;
            rom[29364] = 8'h04 ;
            rom[29365] = 8'hf5 ;
            rom[29366] = 8'h02 ;
            rom[29367] = 8'hd4 ;
            rom[29368] = 8'h15 ;
            rom[29369] = 8'h06 ;
            rom[29370] = 8'heb ;
            rom[29371] = 8'h14 ;
            rom[29372] = 8'hff ;
            rom[29373] = 8'h07 ;
            rom[29374] = 8'hc2 ;
            rom[29375] = 8'h04 ;
            rom[29376] = 8'h18 ;
            rom[29377] = 8'h04 ;
            rom[29378] = 8'hff ;
            rom[29379] = 8'hfe ;
            rom[29380] = 8'he0 ;
            rom[29381] = 8'he0 ;
            rom[29382] = 8'hfa ;
            rom[29383] = 8'hc7 ;
            rom[29384] = 8'hf8 ;
            rom[29385] = 8'h07 ;
            rom[29386] = 8'hff ;
            rom[29387] = 8'h1e ;
            rom[29388] = 8'h09 ;
            rom[29389] = 8'h1d ;
            rom[29390] = 8'he4 ;
            rom[29391] = 8'h03 ;
            rom[29392] = 8'h03 ;
            rom[29393] = 8'h0f ;
            rom[29394] = 8'hde ;
            rom[29395] = 8'hfe ;
            rom[29396] = 8'h30 ;
            rom[29397] = 8'h01 ;
            rom[29398] = 8'he7 ;
            rom[29399] = 8'ha8 ;
            rom[29400] = 8'h00 ;
            rom[29401] = 8'h02 ;
            rom[29402] = 8'h0b ;
            rom[29403] = 8'hf4 ;
            rom[29404] = 8'h01 ;
            rom[29405] = 8'h14 ;
            rom[29406] = 8'he2 ;
            rom[29407] = 8'he8 ;
            rom[29408] = 8'hff ;
            rom[29409] = 8'hec ;
            rom[29410] = 8'h18 ;
            rom[29411] = 8'h15 ;
            rom[29412] = 8'h06 ;
            rom[29413] = 8'h03 ;
            rom[29414] = 8'h14 ;
            rom[29415] = 8'h06 ;
            rom[29416] = 8'he5 ;
            rom[29417] = 8'hc7 ;
            rom[29418] = 8'hdf ;
            rom[29419] = 8'h1a ;
            rom[29420] = 8'hdd ;
            rom[29421] = 8'h03 ;
            rom[29422] = 8'h0d ;
            rom[29423] = 8'hfc ;
            rom[29424] = 8'h13 ;
            rom[29425] = 8'heb ;
            rom[29426] = 8'h07 ;
            rom[29427] = 8'hf4 ;
            rom[29428] = 8'h13 ;
            rom[29429] = 8'hde ;
            rom[29430] = 8'h00 ;
            rom[29431] = 8'h00 ;
            rom[29432] = 8'hcf ;
            rom[29433] = 8'h06 ;
            rom[29434] = 8'hf9 ;
            rom[29435] = 8'h10 ;
            rom[29436] = 8'hd9 ;
            rom[29437] = 8'hc1 ;
            rom[29438] = 8'hba ;
            rom[29439] = 8'h06 ;
            rom[29440] = 8'h06 ;
            rom[29441] = 8'hdc ;
            rom[29442] = 8'hee ;
            rom[29443] = 8'h03 ;
            rom[29444] = 8'h16 ;
            rom[29445] = 8'hfa ;
            rom[29446] = 8'hcd ;
            rom[29447] = 8'h15 ;
            rom[29448] = 8'hf3 ;
            rom[29449] = 8'he2 ;
            rom[29450] = 8'h06 ;
            rom[29451] = 8'he0 ;
            rom[29452] = 8'h11 ;
            rom[29453] = 8'he3 ;
            rom[29454] = 8'h12 ;
            rom[29455] = 8'h02 ;
            rom[29456] = 8'hc6 ;
            rom[29457] = 8'h07 ;
            rom[29458] = 8'hef ;
            rom[29459] = 8'hf9 ;
            rom[29460] = 8'hfb ;
            rom[29461] = 8'hf1 ;
            rom[29462] = 8'hf3 ;
            rom[29463] = 8'he0 ;
            rom[29464] = 8'h08 ;
            rom[29465] = 8'h03 ;
            rom[29466] = 8'h08 ;
            rom[29467] = 8'hf6 ;
            rom[29468] = 8'hfb ;
            rom[29469] = 8'h02 ;
            rom[29470] = 8'hef ;
            rom[29471] = 8'h23 ;
            rom[29472] = 8'h19 ;
            rom[29473] = 8'hb8 ;
            rom[29474] = 8'hc2 ;
            rom[29475] = 8'h30 ;
            rom[29476] = 8'hf6 ;
            rom[29477] = 8'he5 ;
            rom[29478] = 8'h0a ;
            rom[29479] = 8'h09 ;
            rom[29480] = 8'hf8 ;
            rom[29481] = 8'hf4 ;
            rom[29482] = 8'h22 ;
            rom[29483] = 8'h02 ;
            rom[29484] = 8'hfc ;
            rom[29485] = 8'hdc ;
            rom[29486] = 8'h17 ;
            rom[29487] = 8'h12 ;
            rom[29488] = 8'h09 ;
            rom[29489] = 8'hf9 ;
            rom[29490] = 8'he0 ;
            rom[29491] = 8'h1e ;
            rom[29492] = 8'hfa ;
            rom[29493] = 8'h22 ;
            rom[29494] = 8'h12 ;
            rom[29495] = 8'hdd ;
            rom[29496] = 8'hd2 ;
            rom[29497] = 8'h22 ;
            rom[29498] = 8'hfa ;
            rom[29499] = 8'hff ;
            rom[29500] = 8'hd4 ;
            rom[29501] = 8'hf9 ;
            rom[29502] = 8'he9 ;
            rom[29503] = 8'h05 ;
            rom[29504] = 8'hd0 ;
            rom[29505] = 8'h25 ;
            rom[29506] = 8'hef ;
            rom[29507] = 8'hf4 ;
            rom[29508] = 8'h02 ;
            rom[29509] = 8'hfe ;
            rom[29510] = 8'hdd ;
            rom[29511] = 8'h2e ;
            rom[29512] = 8'h03 ;
            rom[29513] = 8'hee ;
            rom[29514] = 8'hf9 ;
            rom[29515] = 8'hfc ;
            rom[29516] = 8'he0 ;
            rom[29517] = 8'hf0 ;
            rom[29518] = 8'he7 ;
            rom[29519] = 8'h03 ;
            rom[29520] = 8'h15 ;
            rom[29521] = 8'hfd ;
            rom[29522] = 8'h11 ;
            rom[29523] = 8'he3 ;
            rom[29524] = 8'he6 ;
            rom[29525] = 8'h1a ;
            rom[29526] = 8'hf8 ;
            rom[29527] = 8'h0a ;
            rom[29528] = 8'hec ;
            rom[29529] = 8'h03 ;
            rom[29530] = 8'h11 ;
            rom[29531] = 8'h06 ;
            rom[29532] = 8'hf6 ;
            rom[29533] = 8'hdc ;
            rom[29534] = 8'h26 ;
            rom[29535] = 8'hfa ;
            rom[29536] = 8'hcc ;
            rom[29537] = 8'h0d ;
            rom[29538] = 8'hea ;
            rom[29539] = 8'hbe ;
            rom[29540] = 8'h00 ;
            rom[29541] = 8'hcf ;
            rom[29542] = 8'hfe ;
            rom[29543] = 8'h09 ;
            rom[29544] = 8'h18 ;
            rom[29545] = 8'h06 ;
            rom[29546] = 8'he5 ;
            rom[29547] = 8'h1d ;
            rom[29548] = 8'h03 ;
            rom[29549] = 8'h15 ;
            rom[29550] = 8'hf6 ;
            rom[29551] = 8'h1b ;
            rom[29552] = 8'h12 ;
            rom[29553] = 8'h1d ;
            rom[29554] = 8'h0a ;
            rom[29555] = 8'hfa ;
            rom[29556] = 8'h02 ;
            rom[29557] = 8'hf6 ;
            rom[29558] = 8'hf1 ;
            rom[29559] = 8'h22 ;
            rom[29560] = 8'h06 ;
            rom[29561] = 8'h02 ;
            rom[29562] = 8'h0f ;
            rom[29563] = 8'hc3 ;
            rom[29564] = 8'h14 ;
            rom[29565] = 8'hf8 ;
            rom[29566] = 8'hf2 ;
            rom[29567] = 8'he0 ;
            rom[29568] = 8'hf3 ;
            rom[29569] = 8'h08 ;
            rom[29570] = 8'hfe ;
            rom[29571] = 8'hcc ;
            rom[29572] = 8'hbe ;
            rom[29573] = 8'hed ;
            rom[29574] = 8'h01 ;
            rom[29575] = 8'h13 ;
            rom[29576] = 8'hfc ;
            rom[29577] = 8'he6 ;
            rom[29578] = 8'hec ;
            rom[29579] = 8'h07 ;
            rom[29580] = 8'hec ;
            rom[29581] = 8'he8 ;
            rom[29582] = 8'h0b ;
            rom[29583] = 8'he6 ;
            rom[29584] = 8'he0 ;
            rom[29585] = 8'h18 ;
            rom[29586] = 8'hca ;
            rom[29587] = 8'h06 ;
            rom[29588] = 8'h0f ;
            rom[29589] = 8'h2d ;
            rom[29590] = 8'hff ;
            rom[29591] = 8'h11 ;
            rom[29592] = 8'hf8 ;
            rom[29593] = 8'hde ;
            rom[29594] = 8'h12 ;
            rom[29595] = 8'h09 ;
            rom[29596] = 8'h09 ;
            rom[29597] = 8'hf7 ;
            rom[29598] = 8'hf9 ;
            rom[29599] = 8'he4 ;
            rom[29600] = 8'hda ;
            rom[29601] = 8'h05 ;
            rom[29602] = 8'h00 ;
            rom[29603] = 8'h11 ;
            rom[29604] = 8'h37 ;
            rom[29605] = 8'h0f ;
            rom[29606] = 8'h08 ;
            rom[29607] = 8'hbc ;
            rom[29608] = 8'hf0 ;
            rom[29609] = 8'he6 ;
            rom[29610] = 8'hff ;
            rom[29611] = 8'hf6 ;
            rom[29612] = 8'h27 ;
            rom[29613] = 8'hfe ;
            rom[29614] = 8'hee ;
            rom[29615] = 8'he3 ;
            rom[29616] = 8'he2 ;
            rom[29617] = 8'he4 ;
            rom[29618] = 8'hdb ;
            rom[29619] = 8'hde ;
            rom[29620] = 8'hf9 ;
            rom[29621] = 8'hdd ;
            rom[29622] = 8'hed ;
            rom[29623] = 8'h16 ;
            rom[29624] = 8'he7 ;
            rom[29625] = 8'h0d ;
            rom[29626] = 8'hdc ;
            rom[29627] = 8'hfb ;
            rom[29628] = 8'hfd ;
            rom[29629] = 8'hc8 ;
            rom[29630] = 8'he8 ;
            rom[29631] = 8'heb ;
            rom[29632] = 8'hfb ;
            rom[29633] = 8'h04 ;
            rom[29634] = 8'he6 ;
            rom[29635] = 8'he9 ;
            rom[29636] = 8'h07 ;
            rom[29637] = 8'h0c ;
            rom[29638] = 8'hf2 ;
            rom[29639] = 8'h04 ;
            rom[29640] = 8'hfe ;
            rom[29641] = 8'h08 ;
            rom[29642] = 8'h20 ;
            rom[29643] = 8'h02 ;
            rom[29644] = 8'hfc ;
            rom[29645] = 8'h22 ;
            rom[29646] = 8'hf4 ;
            rom[29647] = 8'h08 ;
            rom[29648] = 8'hfb ;
            rom[29649] = 8'h01 ;
            rom[29650] = 8'h04 ;
            rom[29651] = 8'hf1 ;
            rom[29652] = 8'h03 ;
            rom[29653] = 8'hdd ;
            rom[29654] = 8'h02 ;
            rom[29655] = 8'h0c ;
            rom[29656] = 8'he5 ;
            rom[29657] = 8'h0d ;
            rom[29658] = 8'h06 ;
            rom[29659] = 8'hcf ;
            rom[29660] = 8'hf8 ;
            rom[29661] = 8'he8 ;
            rom[29662] = 8'h04 ;
            rom[29663] = 8'hf6 ;
            rom[29664] = 8'he4 ;
            rom[29665] = 8'h15 ;
            rom[29666] = 8'hf8 ;
            rom[29667] = 8'h0a ;
            rom[29668] = 8'hd5 ;
            rom[29669] = 8'hed ;
            rom[29670] = 8'h15 ;
            rom[29671] = 8'h16 ;
            rom[29672] = 8'hed ;
            rom[29673] = 8'h0a ;
            rom[29674] = 8'hda ;
            rom[29675] = 8'h19 ;
            rom[29676] = 8'hdc ;
            rom[29677] = 8'h35 ;
            rom[29678] = 8'h01 ;
            rom[29679] = 8'h14 ;
            rom[29680] = 8'h09 ;
            rom[29681] = 8'h09 ;
            rom[29682] = 8'he5 ;
            rom[29683] = 8'h00 ;
            rom[29684] = 8'h17 ;
            rom[29685] = 8'h2d ;
            rom[29686] = 8'h2c ;
            rom[29687] = 8'heb ;
            rom[29688] = 8'he8 ;
            rom[29689] = 8'h18 ;
            rom[29690] = 8'hd8 ;
            rom[29691] = 8'h04 ;
            rom[29692] = 8'heb ;
            rom[29693] = 8'hf3 ;
            rom[29694] = 8'h18 ;
            rom[29695] = 8'hfe ;
            rom[29696] = 8'h1b ;
            rom[29697] = 8'hfa ;
            rom[29698] = 8'hd6 ;
            rom[29699] = 8'hf9 ;
            rom[29700] = 8'hee ;
            rom[29701] = 8'hfd ;
            rom[29702] = 8'hca ;
            rom[29703] = 8'h05 ;
            rom[29704] = 8'hfb ;
            rom[29705] = 8'hf2 ;
            rom[29706] = 8'h0c ;
            rom[29707] = 8'hea ;
            rom[29708] = 8'hfe ;
            rom[29709] = 8'hf3 ;
            rom[29710] = 8'h0f ;
            rom[29711] = 8'hf9 ;
            rom[29712] = 8'heb ;
            rom[29713] = 8'hec ;
            rom[29714] = 8'h08 ;
            rom[29715] = 8'h0e ;
            rom[29716] = 8'hdb ;
            rom[29717] = 8'heb ;
            rom[29718] = 8'hf2 ;
            rom[29719] = 8'h0b ;
            rom[29720] = 8'h00 ;
            rom[29721] = 8'hf5 ;
            rom[29722] = 8'he1 ;
            rom[29723] = 8'hfd ;
            rom[29724] = 8'h00 ;
            rom[29725] = 8'hfa ;
            rom[29726] = 8'h0f ;
            rom[29727] = 8'he7 ;
            rom[29728] = 8'hee ;
            rom[29729] = 8'h09 ;
            rom[29730] = 8'he5 ;
            rom[29731] = 8'h2d ;
            rom[29732] = 8'he5 ;
            rom[29733] = 8'hce ;
            rom[29734] = 8'hce ;
            rom[29735] = 8'h00 ;
            rom[29736] = 8'hf5 ;
            rom[29737] = 8'h15 ;
            rom[29738] = 8'h10 ;
            rom[29739] = 8'h23 ;
            rom[29740] = 8'hc0 ;
            rom[29741] = 8'h17 ;
            rom[29742] = 8'hb5 ;
            rom[29743] = 8'h2b ;
            rom[29744] = 8'hfc ;
            rom[29745] = 8'h07 ;
            rom[29746] = 8'he5 ;
            rom[29747] = 8'h17 ;
            rom[29748] = 8'hf7 ;
            rom[29749] = 8'hf8 ;
            rom[29750] = 8'h11 ;
            rom[29751] = 8'h0a ;
            rom[29752] = 8'h0f ;
            rom[29753] = 8'he3 ;
            rom[29754] = 8'h19 ;
            rom[29755] = 8'heb ;
            rom[29756] = 8'hf8 ;
            rom[29757] = 8'h25 ;
            rom[29758] = 8'h0e ;
            rom[29759] = 8'hea ;
            rom[29760] = 8'he9 ;
            rom[29761] = 8'hea ;
            rom[29762] = 8'h03 ;
            rom[29763] = 8'h16 ;
            rom[29764] = 8'h0b ;
            rom[29765] = 8'h10 ;
            rom[29766] = 8'he9 ;
            rom[29767] = 8'hef ;
            rom[29768] = 8'hf4 ;
            rom[29769] = 8'h17 ;
            rom[29770] = 8'hdf ;
            rom[29771] = 8'hfb ;
            rom[29772] = 8'he5 ;
            rom[29773] = 8'h09 ;
            rom[29774] = 8'heb ;
            rom[29775] = 8'hcd ;
            rom[29776] = 8'h09 ;
            rom[29777] = 8'hff ;
            rom[29778] = 8'h19 ;
            rom[29779] = 8'hea ;
            rom[29780] = 8'h0a ;
            rom[29781] = 8'h07 ;
            rom[29782] = 8'h06 ;
            rom[29783] = 8'hf9 ;
            rom[29784] = 8'hf8 ;
            rom[29785] = 8'hdf ;
            rom[29786] = 8'hdd ;
            rom[29787] = 8'he9 ;
            rom[29788] = 8'hf9 ;
            rom[29789] = 8'h06 ;
            rom[29790] = 8'h03 ;
            rom[29791] = 8'hcb ;
            rom[29792] = 8'hfa ;
            rom[29793] = 8'h0f ;
            rom[29794] = 8'h00 ;
            rom[29795] = 8'hfb ;
            rom[29796] = 8'hf4 ;
            rom[29797] = 8'hf4 ;
            rom[29798] = 8'hf4 ;
            rom[29799] = 8'hf0 ;
            rom[29800] = 8'he9 ;
            rom[29801] = 8'h11 ;
            rom[29802] = 8'hf2 ;
            rom[29803] = 8'h14 ;
            rom[29804] = 8'hfb ;
            rom[29805] = 8'h0c ;
            rom[29806] = 8'h03 ;
            rom[29807] = 8'hf2 ;
            rom[29808] = 8'hd2 ;
            rom[29809] = 8'hfc ;
            rom[29810] = 8'hde ;
            rom[29811] = 8'h00 ;
            rom[29812] = 8'he9 ;
            rom[29813] = 8'h09 ;
            rom[29814] = 8'he2 ;
            rom[29815] = 8'h0d ;
            rom[29816] = 8'he1 ;
            rom[29817] = 8'hdc ;
            rom[29818] = 8'hea ;
            rom[29819] = 8'h0a ;
            rom[29820] = 8'h00 ;
            rom[29821] = 8'he0 ;
            rom[29822] = 8'hfc ;
            rom[29823] = 8'hf2 ;
            rom[29824] = 8'hf0 ;
            rom[29825] = 8'hf5 ;
            rom[29826] = 8'h0f ;
            rom[29827] = 8'hf9 ;
            rom[29828] = 8'hf6 ;
            rom[29829] = 8'hf3 ;
            rom[29830] = 8'h15 ;
            rom[29831] = 8'hd3 ;
            rom[29832] = 8'hc7 ;
            rom[29833] = 8'h0e ;
            rom[29834] = 8'hee ;
            rom[29835] = 8'h09 ;
            rom[29836] = 8'hdc ;
            rom[29837] = 8'h1d ;
            rom[29838] = 8'hf7 ;
            rom[29839] = 8'h04 ;
            rom[29840] = 8'h09 ;
            rom[29841] = 8'h23 ;
            rom[29842] = 8'hac ;
            rom[29843] = 8'hcc ;
            rom[29844] = 8'h2d ;
            rom[29845] = 8'h1a ;
            rom[29846] = 8'h02 ;
            rom[29847] = 8'hfa ;
            rom[29848] = 8'h15 ;
            rom[29849] = 8'h09 ;
            rom[29850] = 8'hfe ;
            rom[29851] = 8'hf8 ;
            rom[29852] = 8'heb ;
            rom[29853] = 8'hf9 ;
            rom[29854] = 8'hfb ;
            rom[29855] = 8'he4 ;
            rom[29856] = 8'he6 ;
            rom[29857] = 8'h10 ;
            rom[29858] = 8'hde ;
            rom[29859] = 8'h12 ;
            rom[29860] = 8'h2b ;
            rom[29861] = 8'he7 ;
            rom[29862] = 8'h18 ;
            rom[29863] = 8'hf0 ;
            rom[29864] = 8'h21 ;
            rom[29865] = 8'hfa ;
            rom[29866] = 8'h00 ;
            rom[29867] = 8'he7 ;
            rom[29868] = 8'h02 ;
            rom[29869] = 8'hf4 ;
            rom[29870] = 8'hfd ;
            rom[29871] = 8'hc0 ;
            rom[29872] = 8'hd9 ;
            rom[29873] = 8'he8 ;
            rom[29874] = 8'hcb ;
            rom[29875] = 8'heb ;
            rom[29876] = 8'h09 ;
            rom[29877] = 8'hba ;
            rom[29878] = 8'hee ;
            rom[29879] = 8'hf0 ;
            rom[29880] = 8'h0b ;
            rom[29881] = 8'hf8 ;
            rom[29882] = 8'hde ;
            rom[29883] = 8'h03 ;
            rom[29884] = 8'h01 ;
            rom[29885] = 8'hcd ;
            rom[29886] = 8'hf9 ;
            rom[29887] = 8'h03 ;
            rom[29888] = 8'hf7 ;
            rom[29889] = 8'h26 ;
            rom[29890] = 8'h10 ;
            rom[29891] = 8'h0c ;
            rom[29892] = 8'h15 ;
            rom[29893] = 8'hfb ;
            rom[29894] = 8'hc6 ;
            rom[29895] = 8'hf2 ;
            rom[29896] = 8'hf3 ;
            rom[29897] = 8'hed ;
            rom[29898] = 8'h21 ;
            rom[29899] = 8'h0b ;
            rom[29900] = 8'h07 ;
            rom[29901] = 8'h03 ;
            rom[29902] = 8'h0e ;
            rom[29903] = 8'h0c ;
            rom[29904] = 8'he1 ;
            rom[29905] = 8'h02 ;
            rom[29906] = 8'hcf ;
            rom[29907] = 8'h0c ;
            rom[29908] = 8'hf1 ;
            rom[29909] = 8'hf2 ;
            rom[29910] = 8'hf9 ;
            rom[29911] = 8'h0a ;
            rom[29912] = 8'h1d ;
            rom[29913] = 8'hf4 ;
            rom[29914] = 8'hf9 ;
            rom[29915] = 8'hef ;
            rom[29916] = 8'h13 ;
            rom[29917] = 8'h0f ;
            rom[29918] = 8'h12 ;
            rom[29919] = 8'hff ;
            rom[29920] = 8'he7 ;
            rom[29921] = 8'hef ;
            rom[29922] = 8'hcc ;
            rom[29923] = 8'he7 ;
            rom[29924] = 8'h05 ;
            rom[29925] = 8'hf6 ;
            rom[29926] = 8'he0 ;
            rom[29927] = 8'h19 ;
            rom[29928] = 8'hd6 ;
            rom[29929] = 8'hf2 ;
            rom[29930] = 8'hee ;
            rom[29931] = 8'he0 ;
            rom[29932] = 8'he3 ;
            rom[29933] = 8'he3 ;
            rom[29934] = 8'h05 ;
            rom[29935] = 8'hfa ;
            rom[29936] = 8'h20 ;
            rom[29937] = 8'h18 ;
            rom[29938] = 8'h0f ;
            rom[29939] = 8'hfe ;
            rom[29940] = 8'h17 ;
            rom[29941] = 8'h0b ;
            rom[29942] = 8'h11 ;
            rom[29943] = 8'h05 ;
            rom[29944] = 8'h04 ;
            rom[29945] = 8'h0b ;
            rom[29946] = 8'h23 ;
            rom[29947] = 8'hce ;
            rom[29948] = 8'hed ;
            rom[29949] = 8'h17 ;
            rom[29950] = 8'hd1 ;
            rom[29951] = 8'hbc ;
            rom[29952] = 8'hcc ;
            rom[29953] = 8'he2 ;
            rom[29954] = 8'he6 ;
            rom[29955] = 8'h09 ;
            rom[29956] = 8'hf0 ;
            rom[29957] = 8'h0a ;
            rom[29958] = 8'hf0 ;
            rom[29959] = 8'h16 ;
            rom[29960] = 8'hee ;
            rom[29961] = 8'h1d ;
            rom[29962] = 8'hf2 ;
            rom[29963] = 8'h04 ;
            rom[29964] = 8'h0c ;
            rom[29965] = 8'hd8 ;
            rom[29966] = 8'hf9 ;
            rom[29967] = 8'h07 ;
            rom[29968] = 8'h1c ;
            rom[29969] = 8'hf1 ;
            rom[29970] = 8'h02 ;
            rom[29971] = 8'h1c ;
            rom[29972] = 8'h13 ;
            rom[29973] = 8'he1 ;
            rom[29974] = 8'hf8 ;
            rom[29975] = 8'h2a ;
            rom[29976] = 8'hfa ;
            rom[29977] = 8'h0c ;
            rom[29978] = 8'hfc ;
            rom[29979] = 8'h06 ;
            rom[29980] = 8'hdb ;
            rom[29981] = 8'h0a ;
            rom[29982] = 8'hfb ;
            rom[29983] = 8'hfd ;
            rom[29984] = 8'hf4 ;
            rom[29985] = 8'hf3 ;
            rom[29986] = 8'h02 ;
            rom[29987] = 8'hed ;
            rom[29988] = 8'he8 ;
            rom[29989] = 8'hed ;
            rom[29990] = 8'he8 ;
            rom[29991] = 8'h0a ;
            rom[29992] = 8'h04 ;
            rom[29993] = 8'he6 ;
            rom[29994] = 8'hfe ;
            rom[29995] = 8'h12 ;
            rom[29996] = 8'hee ;
            rom[29997] = 8'he5 ;
            rom[29998] = 8'h09 ;
            rom[29999] = 8'hfa ;
            rom[30000] = 8'h0d ;
            rom[30001] = 8'hd9 ;
            rom[30002] = 8'h06 ;
            rom[30003] = 8'h04 ;
            rom[30004] = 8'hed ;
            rom[30005] = 8'h1d ;
            rom[30006] = 8'h18 ;
            rom[30007] = 8'hef ;
            rom[30008] = 8'hf1 ;
            rom[30009] = 8'h13 ;
            rom[30010] = 8'h08 ;
            rom[30011] = 8'h01 ;
            rom[30012] = 8'hfb ;
            rom[30013] = 8'hff ;
            rom[30014] = 8'hf3 ;
            rom[30015] = 8'hf3 ;
            rom[30016] = 8'heb ;
            rom[30017] = 8'hda ;
            rom[30018] = 8'he5 ;
            rom[30019] = 8'hfe ;
            rom[30020] = 8'hf0 ;
            rom[30021] = 8'he7 ;
            rom[30022] = 8'h0d ;
            rom[30023] = 8'hff ;
            rom[30024] = 8'hf8 ;
            rom[30025] = 8'hf1 ;
            rom[30026] = 8'h20 ;
            rom[30027] = 8'h1e ;
            rom[30028] = 8'hf5 ;
            rom[30029] = 8'heb ;
            rom[30030] = 8'hcb ;
            rom[30031] = 8'hdf ;
            rom[30032] = 8'hfb ;
            rom[30033] = 8'hfc ;
            rom[30034] = 8'hf9 ;
            rom[30035] = 8'hf5 ;
            rom[30036] = 8'h0b ;
            rom[30037] = 8'h02 ;
            rom[30038] = 8'h2e ;
            rom[30039] = 8'he9 ;
            rom[30040] = 8'hf0 ;
            rom[30041] = 8'h1e ;
            rom[30042] = 8'h0d ;
            rom[30043] = 8'hf5 ;
            rom[30044] = 8'hfa ;
            rom[30045] = 8'h06 ;
            rom[30046] = 8'h18 ;
            rom[30047] = 8'hf6 ;
            rom[30048] = 8'h1e ;
            rom[30049] = 8'hf8 ;
            rom[30050] = 8'hf0 ;
            rom[30051] = 8'he1 ;
            rom[30052] = 8'he2 ;
            rom[30053] = 8'h19 ;
            rom[30054] = 8'h0a ;
            rom[30055] = 8'he5 ;
            rom[30056] = 8'h01 ;
            rom[30057] = 8'hb7 ;
            rom[30058] = 8'heb ;
            rom[30059] = 8'h14 ;
            rom[30060] = 8'hec ;
            rom[30061] = 8'he9 ;
            rom[30062] = 8'hf2 ;
            rom[30063] = 8'hcc ;
            rom[30064] = 8'hfb ;
            rom[30065] = 8'hd7 ;
            rom[30066] = 8'h02 ;
            rom[30067] = 8'hcd ;
            rom[30068] = 8'h04 ;
            rom[30069] = 8'hc0 ;
            rom[30070] = 8'hf2 ;
            rom[30071] = 8'hf3 ;
            rom[30072] = 8'hed ;
            rom[30073] = 8'hfe ;
            rom[30074] = 8'hfc ;
            rom[30075] = 8'hff ;
            rom[30076] = 8'hd8 ;
            rom[30077] = 8'hea ;
            rom[30078] = 8'heb ;
            rom[30079] = 8'h1b ;
            rom[30080] = 8'hef ;
            rom[30081] = 8'h08 ;
            rom[30082] = 8'hff ;
            rom[30083] = 8'hfc ;
            rom[30084] = 8'h07 ;
            rom[30085] = 8'heb ;
            rom[30086] = 8'h1d ;
            rom[30087] = 8'hed ;
            rom[30088] = 8'he5 ;
            rom[30089] = 8'hff ;
            rom[30090] = 8'hf2 ;
            rom[30091] = 8'he7 ;
            rom[30092] = 8'he7 ;
            rom[30093] = 8'h09 ;
            rom[30094] = 8'h1b ;
            rom[30095] = 8'hef ;
            rom[30096] = 8'hf4 ;
            rom[30097] = 8'had ;
            rom[30098] = 8'hff ;
            rom[30099] = 8'h16 ;
            rom[30100] = 8'h0e ;
            rom[30101] = 8'h07 ;
            rom[30102] = 8'hf2 ;
            rom[30103] = 8'heb ;
            rom[30104] = 8'hfb ;
            rom[30105] = 8'h1c ;
            rom[30106] = 8'hfe ;
            rom[30107] = 8'hda ;
            rom[30108] = 8'heb ;
            rom[30109] = 8'h04 ;
            rom[30110] = 8'h08 ;
            rom[30111] = 8'hd1 ;
            rom[30112] = 8'h0a ;
            rom[30113] = 8'hfb ;
            rom[30114] = 8'hfa ;
            rom[30115] = 8'hdf ;
            rom[30116] = 8'h1b ;
            rom[30117] = 8'hec ;
            rom[30118] = 8'hec ;
            rom[30119] = 8'h0c ;
            rom[30120] = 8'hf1 ;
            rom[30121] = 8'hf0 ;
            rom[30122] = 8'h06 ;
            rom[30123] = 8'hfa ;
            rom[30124] = 8'he1 ;
            rom[30125] = 8'h06 ;
            rom[30126] = 8'hfa ;
            rom[30127] = 8'he8 ;
            rom[30128] = 8'hd9 ;
            rom[30129] = 8'h08 ;
            rom[30130] = 8'h0c ;
            rom[30131] = 8'he3 ;
            rom[30132] = 8'hf7 ;
            rom[30133] = 8'hea ;
            rom[30134] = 8'he2 ;
            rom[30135] = 8'hf4 ;
            rom[30136] = 8'hf6 ;
            rom[30137] = 8'h1e ;
            rom[30138] = 8'heb ;
            rom[30139] = 8'hf5 ;
            rom[30140] = 8'hf3 ;
            rom[30141] = 8'he0 ;
            rom[30142] = 8'hc9 ;
            rom[30143] = 8'he2 ;
            rom[30144] = 8'hef ;
            rom[30145] = 8'hf1 ;
            rom[30146] = 8'h08 ;
            rom[30147] = 8'hf5 ;
            rom[30148] = 8'hf2 ;
            rom[30149] = 8'hf3 ;
            rom[30150] = 8'hfa ;
            rom[30151] = 8'hf4 ;
            rom[30152] = 8'h03 ;
            rom[30153] = 8'he9 ;
            rom[30154] = 8'hf2 ;
            rom[30155] = 8'he9 ;
            rom[30156] = 8'he6 ;
            rom[30157] = 8'h04 ;
            rom[30158] = 8'hdc ;
            rom[30159] = 8'he1 ;
            rom[30160] = 8'hfa ;
            rom[30161] = 8'he8 ;
            rom[30162] = 8'he0 ;
            rom[30163] = 8'h17 ;
            rom[30164] = 8'he0 ;
            rom[30165] = 8'hf4 ;
            rom[30166] = 8'hfe ;
            rom[30167] = 8'hed ;
            rom[30168] = 8'heb ;
            rom[30169] = 8'he3 ;
            rom[30170] = 8'hd9 ;
            rom[30171] = 8'hdc ;
            rom[30172] = 8'he8 ;
            rom[30173] = 8'hfa ;
            rom[30174] = 8'he2 ;
            rom[30175] = 8'hd3 ;
            rom[30176] = 8'h10 ;
            rom[30177] = 8'h07 ;
            rom[30178] = 8'he1 ;
            rom[30179] = 8'h09 ;
            rom[30180] = 8'h06 ;
            rom[30181] = 8'h10 ;
            rom[30182] = 8'hf4 ;
            rom[30183] = 8'hde ;
            rom[30184] = 8'he8 ;
            rom[30185] = 8'hec ;
            rom[30186] = 8'h19 ;
            rom[30187] = 8'h14 ;
            rom[30188] = 8'hdb ;
            rom[30189] = 8'h06 ;
            rom[30190] = 8'hf6 ;
            rom[30191] = 8'hf8 ;
            rom[30192] = 8'h01 ;
            rom[30193] = 8'hbb ;
            rom[30194] = 8'h10 ;
            rom[30195] = 8'hf4 ;
            rom[30196] = 8'hd0 ;
            rom[30197] = 8'hfd ;
            rom[30198] = 8'hb0 ;
            rom[30199] = 8'hd1 ;
            rom[30200] = 8'he5 ;
            rom[30201] = 8'hdf ;
            rom[30202] = 8'h12 ;
            rom[30203] = 8'hec ;
            rom[30204] = 8'hc5 ;
            rom[30205] = 8'hb0 ;
            rom[30206] = 8'h06 ;
            rom[30207] = 8'h01 ;
            rom[30208] = 8'hd6 ;
            rom[30209] = 8'hb6 ;
            rom[30210] = 8'hd4 ;
            rom[30211] = 8'h05 ;
            rom[30212] = 8'hed ;
            rom[30213] = 8'h03 ;
            rom[30214] = 8'h12 ;
            rom[30215] = 8'h09 ;
            rom[30216] = 8'he9 ;
            rom[30217] = 8'hdc ;
            rom[30218] = 8'he5 ;
            rom[30219] = 8'he8 ;
            rom[30220] = 8'he5 ;
            rom[30221] = 8'h12 ;
            rom[30222] = 8'h1f ;
            rom[30223] = 8'hcd ;
            rom[30224] = 8'hf3 ;
            rom[30225] = 8'h10 ;
            rom[30226] = 8'hd8 ;
            rom[30227] = 8'had ;
            rom[30228] = 8'hea ;
            rom[30229] = 8'he7 ;
            rom[30230] = 8'h02 ;
            rom[30231] = 8'he2 ;
            rom[30232] = 8'h1f ;
            rom[30233] = 8'hf1 ;
            rom[30234] = 8'h0f ;
            rom[30235] = 8'hfa ;
            rom[30236] = 8'h19 ;
            rom[30237] = 8'h00 ;
            rom[30238] = 8'hf6 ;
            rom[30239] = 8'h09 ;
            rom[30240] = 8'h07 ;
            rom[30241] = 8'h0d ;
            rom[30242] = 8'hde ;
            rom[30243] = 8'hcf ;
            rom[30244] = 8'hfc ;
            rom[30245] = 8'hf1 ;
            rom[30246] = 8'h16 ;
            rom[30247] = 8'hd3 ;
            rom[30248] = 8'hec ;
            rom[30249] = 8'hf9 ;
            rom[30250] = 8'h05 ;
            rom[30251] = 8'hb8 ;
            rom[30252] = 8'h39 ;
            rom[30253] = 8'h08 ;
            rom[30254] = 8'he2 ;
            rom[30255] = 8'h14 ;
            rom[30256] = 8'hf0 ;
            rom[30257] = 8'hf4 ;
            rom[30258] = 8'h02 ;
            rom[30259] = 8'hfa ;
            rom[30260] = 8'h05 ;
            rom[30261] = 8'h01 ;
            rom[30262] = 8'hd5 ;
            rom[30263] = 8'h28 ;
            rom[30264] = 8'he9 ;
            rom[30265] = 8'hfd ;
            rom[30266] = 8'hc5 ;
            rom[30267] = 8'hc4 ;
            rom[30268] = 8'he4 ;
            rom[30269] = 8'h14 ;
            rom[30270] = 8'hee ;
            rom[30271] = 8'hee ;
            rom[30272] = 8'h23 ;
            rom[30273] = 8'h28 ;
            rom[30274] = 8'h3e ;
            rom[30275] = 8'hdf ;
            rom[30276] = 8'h17 ;
            rom[30277] = 8'he0 ;
            rom[30278] = 8'h0e ;
            rom[30279] = 8'h03 ;
            rom[30280] = 8'hfc ;
            rom[30281] = 8'hea ;
            rom[30282] = 8'h1b ;
            rom[30283] = 8'hf9 ;
            rom[30284] = 8'hc9 ;
            rom[30285] = 8'hf7 ;
            rom[30286] = 8'hf9 ;
            rom[30287] = 8'hfe ;
            rom[30288] = 8'hd6 ;
            rom[30289] = 8'he4 ;
            rom[30290] = 8'he3 ;
            rom[30291] = 8'hfb ;
            rom[30292] = 8'hca ;
            rom[30293] = 8'h04 ;
            rom[30294] = 8'h02 ;
            rom[30295] = 8'h22 ;
            rom[30296] = 8'hf6 ;
            rom[30297] = 8'hf8 ;
            rom[30298] = 8'hdd ;
            rom[30299] = 8'h27 ;
            rom[30300] = 8'hef ;
            rom[30301] = 8'hfe ;
            rom[30302] = 8'he5 ;
            rom[30303] = 8'h08 ;
            rom[30304] = 8'hdc ;
            rom[30305] = 8'hfd ;
            rom[30306] = 8'hcc ;
            rom[30307] = 8'h02 ;
            rom[30308] = 8'hc1 ;
            rom[30309] = 8'hee ;
            rom[30310] = 8'he5 ;
            rom[30311] = 8'hff ;
            rom[30312] = 8'h0c ;
            rom[30313] = 8'hfe ;
            rom[30314] = 8'h0e ;
            rom[30315] = 8'hef ;
            rom[30316] = 8'hfa ;
            rom[30317] = 8'he1 ;
            rom[30318] = 8'hf6 ;
            rom[30319] = 8'h11 ;
            rom[30320] = 8'h06 ;
            rom[30321] = 8'h17 ;
            rom[30322] = 8'h14 ;
            rom[30323] = 8'h12 ;
            rom[30324] = 8'hf1 ;
            rom[30325] = 8'he7 ;
            rom[30326] = 8'h1b ;
            rom[30327] = 8'hf5 ;
            rom[30328] = 8'h02 ;
            rom[30329] = 8'hc3 ;
            rom[30330] = 8'hf7 ;
            rom[30331] = 8'h14 ;
            rom[30332] = 8'h0c ;
            rom[30333] = 8'h27 ;
            rom[30334] = 8'hd9 ;
            rom[30335] = 8'hd8 ;
            rom[30336] = 8'h05 ;
            rom[30337] = 8'he6 ;
            rom[30338] = 8'ha9 ;
            rom[30339] = 8'h1a ;
            rom[30340] = 8'h13 ;
            rom[30341] = 8'hd9 ;
            rom[30342] = 8'h05 ;
            rom[30343] = 8'h29 ;
            rom[30344] = 8'hf0 ;
            rom[30345] = 8'hcf ;
            rom[30346] = 8'hf4 ;
            rom[30347] = 8'h01 ;
            rom[30348] = 8'hdf ;
            rom[30349] = 8'hf4 ;
            rom[30350] = 8'h03 ;
            rom[30351] = 8'h0a ;
            rom[30352] = 8'hf6 ;
            rom[30353] = 8'he8 ;
            rom[30354] = 8'h0f ;
            rom[30355] = 8'hf5 ;
            rom[30356] = 8'he1 ;
            rom[30357] = 8'hfc ;
            rom[30358] = 8'hea ;
            rom[30359] = 8'h2c ;
            rom[30360] = 8'h19 ;
            rom[30361] = 8'hfd ;
            rom[30362] = 8'h0a ;
            rom[30363] = 8'h17 ;
            rom[30364] = 8'he8 ;
            rom[30365] = 8'h1b ;
            rom[30366] = 8'h04 ;
            rom[30367] = 8'hf1 ;
            rom[30368] = 8'h02 ;
            rom[30369] = 8'h1a ;
            rom[30370] = 8'h0e ;
            rom[30371] = 8'hd5 ;
            rom[30372] = 8'he8 ;
            rom[30373] = 8'h0b ;
            rom[30374] = 8'h0b ;
            rom[30375] = 8'hfd ;
            rom[30376] = 8'hec ;
            rom[30377] = 8'h05 ;
            rom[30378] = 8'h20 ;
            rom[30379] = 8'h0d ;
            rom[30380] = 8'hdb ;
            rom[30381] = 8'h0e ;
            rom[30382] = 8'hf7 ;
            rom[30383] = 8'h08 ;
            rom[30384] = 8'hf9 ;
            rom[30385] = 8'h18 ;
            rom[30386] = 8'h00 ;
            rom[30387] = 8'hef ;
            rom[30388] = 8'hfb ;
            rom[30389] = 8'he3 ;
            rom[30390] = 8'hfe ;
            rom[30391] = 8'h1e ;
            rom[30392] = 8'hf8 ;
            rom[30393] = 8'h1a ;
            rom[30394] = 8'he3 ;
            rom[30395] = 8'he8 ;
            rom[30396] = 8'h00 ;
            rom[30397] = 8'h04 ;
            rom[30398] = 8'hf6 ;
            rom[30399] = 8'hc4 ;
            rom[30400] = 8'h11 ;
            rom[30401] = 8'h0a ;
            rom[30402] = 8'hfc ;
            rom[30403] = 8'h06 ;
            rom[30404] = 8'hf7 ;
            rom[30405] = 8'h05 ;
            rom[30406] = 8'hfc ;
            rom[30407] = 8'hf1 ;
            rom[30408] = 8'hff ;
            rom[30409] = 8'h12 ;
            rom[30410] = 8'hf4 ;
            rom[30411] = 8'hf4 ;
            rom[30412] = 8'he3 ;
            rom[30413] = 8'h0e ;
            rom[30414] = 8'he2 ;
            rom[30415] = 8'he7 ;
            rom[30416] = 8'hf6 ;
            rom[30417] = 8'h23 ;
            rom[30418] = 8'hf8 ;
            rom[30419] = 8'h0b ;
            rom[30420] = 8'heb ;
            rom[30421] = 8'hd4 ;
            rom[30422] = 8'h00 ;
            rom[30423] = 8'h3d ;
            rom[30424] = 8'he9 ;
            rom[30425] = 8'h2c ;
            rom[30426] = 8'hd9 ;
            rom[30427] = 8'hdc ;
            rom[30428] = 8'he9 ;
            rom[30429] = 8'he1 ;
            rom[30430] = 8'hf1 ;
            rom[30431] = 8'hfc ;
            rom[30432] = 8'h0f ;
            rom[30433] = 8'h17 ;
            rom[30434] = 8'hce ;
            rom[30435] = 8'h0d ;
            rom[30436] = 8'h17 ;
            rom[30437] = 8'hf1 ;
            rom[30438] = 8'hea ;
            rom[30439] = 8'hba ;
            rom[30440] = 8'h1d ;
            rom[30441] = 8'hd1 ;
            rom[30442] = 8'hd3 ;
            rom[30443] = 8'h01 ;
            rom[30444] = 8'hef ;
            rom[30445] = 8'hdb ;
            rom[30446] = 8'hfb ;
            rom[30447] = 8'hf9 ;
            rom[30448] = 8'hfa ;
            rom[30449] = 8'hd9 ;
            rom[30450] = 8'he7 ;
            rom[30451] = 8'h16 ;
            rom[30452] = 8'hcb ;
            rom[30453] = 8'hf8 ;
            rom[30454] = 8'hdd ;
            rom[30455] = 8'hbf ;
            rom[30456] = 8'h07 ;
            rom[30457] = 8'he9 ;
            rom[30458] = 8'hf9 ;
            rom[30459] = 8'h12 ;
            rom[30460] = 8'hf3 ;
            rom[30461] = 8'hfd ;
            rom[30462] = 8'hfa ;
            rom[30463] = 8'h0d ;
            rom[30464] = 8'h0d ;
            rom[30465] = 8'h1a ;
            rom[30466] = 8'hea ;
            rom[30467] = 8'hdc ;
            rom[30468] = 8'h1e ;
            rom[30469] = 8'hf3 ;
            rom[30470] = 8'hda ;
            rom[30471] = 8'hf7 ;
            rom[30472] = 8'h1d ;
            rom[30473] = 8'he9 ;
            rom[30474] = 8'h16 ;
            rom[30475] = 8'hf3 ;
            rom[30476] = 8'he0 ;
            rom[30477] = 8'h11 ;
            rom[30478] = 8'hfd ;
            rom[30479] = 8'h05 ;
            rom[30480] = 8'heb ;
            rom[30481] = 8'h0a ;
            rom[30482] = 8'h20 ;
            rom[30483] = 8'he7 ;
            rom[30484] = 8'hed ;
            rom[30485] = 8'h08 ;
            rom[30486] = 8'hfd ;
            rom[30487] = 8'h02 ;
            rom[30488] = 8'hb4 ;
            rom[30489] = 8'he4 ;
            rom[30490] = 8'h05 ;
            rom[30491] = 8'hbf ;
            rom[30492] = 8'he0 ;
            rom[30493] = 8'h02 ;
            rom[30494] = 8'hf9 ;
            rom[30495] = 8'h1d ;
            rom[30496] = 8'h28 ;
            rom[30497] = 8'he9 ;
            rom[30498] = 8'h24 ;
            rom[30499] = 8'h1f ;
            rom[30500] = 8'hfa ;
            rom[30501] = 8'he0 ;
            rom[30502] = 8'h11 ;
            rom[30503] = 8'h00 ;
            rom[30504] = 8'h1b ;
            rom[30505] = 8'hf5 ;
            rom[30506] = 8'he3 ;
            rom[30507] = 8'h20 ;
            rom[30508] = 8'hf2 ;
            rom[30509] = 8'hf1 ;
            rom[30510] = 8'h12 ;
            rom[30511] = 8'hf7 ;
            rom[30512] = 8'hfb ;
            rom[30513] = 8'he7 ;
            rom[30514] = 8'he1 ;
            rom[30515] = 8'hf9 ;
            rom[30516] = 8'hf4 ;
            rom[30517] = 8'h01 ;
            rom[30518] = 8'h07 ;
            rom[30519] = 8'h23 ;
            rom[30520] = 8'h09 ;
            rom[30521] = 8'hdc ;
            rom[30522] = 8'hf5 ;
            rom[30523] = 8'hed ;
            rom[30524] = 8'h09 ;
            rom[30525] = 8'he1 ;
            rom[30526] = 8'h08 ;
            rom[30527] = 8'h26 ;
            rom[30528] = 8'hec ;
            rom[30529] = 8'hd5 ;
            rom[30530] = 8'hec ;
            rom[30531] = 8'h15 ;
            rom[30532] = 8'hf3 ;
            rom[30533] = 8'h16 ;
            rom[30534] = 8'hdd ;
            rom[30535] = 8'h1a ;
            rom[30536] = 8'he6 ;
            rom[30537] = 8'hff ;
            rom[30538] = 8'hef ;
            rom[30539] = 8'hf3 ;
            rom[30540] = 8'hfa ;
            rom[30541] = 8'he2 ;
            rom[30542] = 8'hf5 ;
            rom[30543] = 8'heb ;
            rom[30544] = 8'hed ;
            rom[30545] = 8'h04 ;
            rom[30546] = 8'h1a ;
            rom[30547] = 8'he6 ;
            rom[30548] = 8'h1e ;
            rom[30549] = 8'h01 ;
            rom[30550] = 8'hdd ;
            rom[30551] = 8'hfe ;
            rom[30552] = 8'hdd ;
            rom[30553] = 8'h01 ;
            rom[30554] = 8'h17 ;
            rom[30555] = 8'hf8 ;
            rom[30556] = 8'he5 ;
            rom[30557] = 8'h11 ;
            rom[30558] = 8'h0e ;
            rom[30559] = 8'h12 ;
            rom[30560] = 8'hf8 ;
            rom[30561] = 8'h05 ;
            rom[30562] = 8'he8 ;
            rom[30563] = 8'he1 ;
            rom[30564] = 8'hfe ;
            rom[30565] = 8'hfe ;
            rom[30566] = 8'hf8 ;
            rom[30567] = 8'hff ;
            rom[30568] = 8'hec ;
            rom[30569] = 8'h09 ;
            rom[30570] = 8'hee ;
            rom[30571] = 8'hd7 ;
            rom[30572] = 8'h08 ;
            rom[30573] = 8'h00 ;
            rom[30574] = 8'h06 ;
            rom[30575] = 8'hed ;
            rom[30576] = 8'hd4 ;
            rom[30577] = 8'he7 ;
            rom[30578] = 8'h13 ;
            rom[30579] = 8'hf1 ;
            rom[30580] = 8'hfb ;
            rom[30581] = 8'h17 ;
            rom[30582] = 8'heb ;
            rom[30583] = 8'hf2 ;
            rom[30584] = 8'hfe ;
            rom[30585] = 8'he0 ;
            rom[30586] = 8'hf2 ;
            rom[30587] = 8'h09 ;
            rom[30588] = 8'hfc ;
            rom[30589] = 8'hdb ;
            rom[30590] = 8'h11 ;
            rom[30591] = 8'h05 ;
            rom[30592] = 8'h2d ;
            rom[30593] = 8'hf7 ;
            rom[30594] = 8'hf4 ;
            rom[30595] = 8'hfa ;
            rom[30596] = 8'he1 ;
            rom[30597] = 8'hf1 ;
            rom[30598] = 8'h1c ;
            rom[30599] = 8'h31 ;
            rom[30600] = 8'hd2 ;
            rom[30601] = 8'h10 ;
            rom[30602] = 8'he0 ;
            rom[30603] = 8'hf7 ;
            rom[30604] = 8'hf9 ;
            rom[30605] = 8'hd7 ;
            rom[30606] = 8'h08 ;
            rom[30607] = 8'hd3 ;
            rom[30608] = 8'hf2 ;
            rom[30609] = 8'h1f ;
            rom[30610] = 8'h08 ;
            rom[30611] = 8'h0f ;
            rom[30612] = 8'h0d ;
            rom[30613] = 8'hd2 ;
            rom[30614] = 8'heb ;
            rom[30615] = 8'hf0 ;
            rom[30616] = 8'h17 ;
            rom[30617] = 8'h05 ;
            rom[30618] = 8'hf1 ;
            rom[30619] = 8'h06 ;
            rom[30620] = 8'h10 ;
            rom[30621] = 8'hf9 ;
            rom[30622] = 8'h06 ;
            rom[30623] = 8'hf9 ;
            rom[30624] = 8'h13 ;
            rom[30625] = 8'h1d ;
            rom[30626] = 8'h18 ;
            rom[30627] = 8'h14 ;
            rom[30628] = 8'hee ;
            rom[30629] = 8'h04 ;
            rom[30630] = 8'h0c ;
            rom[30631] = 8'hfb ;
            rom[30632] = 8'he7 ;
            rom[30633] = 8'hc1 ;
            rom[30634] = 8'hdf ;
            rom[30635] = 8'hf2 ;
            rom[30636] = 8'hfe ;
            rom[30637] = 8'hfa ;
            rom[30638] = 8'he8 ;
            rom[30639] = 8'h1e ;
            rom[30640] = 8'hfc ;
            rom[30641] = 8'he2 ;
            rom[30642] = 8'h0b ;
            rom[30643] = 8'h0b ;
            rom[30644] = 8'heb ;
            rom[30645] = 8'h21 ;
            rom[30646] = 8'hf6 ;
            rom[30647] = 8'h0c ;
            rom[30648] = 8'hea ;
            rom[30649] = 8'hc9 ;
            rom[30650] = 8'h0b ;
            rom[30651] = 8'h02 ;
            rom[30652] = 8'hd0 ;
            rom[30653] = 8'hfe ;
            rom[30654] = 8'he0 ;
            rom[30655] = 8'h18 ;
            rom[30656] = 8'h13 ;
            rom[30657] = 8'he7 ;
            rom[30658] = 8'h03 ;
            rom[30659] = 8'he3 ;
            rom[30660] = 8'hfb ;
            rom[30661] = 8'hf1 ;
            rom[30662] = 8'hf3 ;
            rom[30663] = 8'hfe ;
            rom[30664] = 8'hf7 ;
            rom[30665] = 8'hf8 ;
            rom[30666] = 8'h0d ;
            rom[30667] = 8'h13 ;
            rom[30668] = 8'hfe ;
            rom[30669] = 8'hf0 ;
            rom[30670] = 8'hed ;
            rom[30671] = 8'hf8 ;
            rom[30672] = 8'h12 ;
            rom[30673] = 8'hec ;
            rom[30674] = 8'h0f ;
            rom[30675] = 8'he4 ;
            rom[30676] = 8'h03 ;
            rom[30677] = 8'h11 ;
            rom[30678] = 8'ha2 ;
            rom[30679] = 8'h05 ;
            rom[30680] = 8'hf6 ;
            rom[30681] = 8'hd6 ;
            rom[30682] = 8'h10 ;
            rom[30683] = 8'h1b ;
            rom[30684] = 8'h04 ;
            rom[30685] = 8'he6 ;
            rom[30686] = 8'h12 ;
            rom[30687] = 8'hf6 ;
            rom[30688] = 8'hec ;
            rom[30689] = 8'hf3 ;
            rom[30690] = 8'h0c ;
            rom[30691] = 8'hf7 ;
            rom[30692] = 8'hd4 ;
            rom[30693] = 8'hff ;
            rom[30694] = 8'h03 ;
            rom[30695] = 8'hfb ;
            rom[30696] = 8'h17 ;
            rom[30697] = 8'h02 ;
            rom[30698] = 8'h17 ;
            rom[30699] = 8'hec ;
            rom[30700] = 8'hff ;
            rom[30701] = 8'h0d ;
            rom[30702] = 8'he9 ;
            rom[30703] = 8'h06 ;
            rom[30704] = 8'h02 ;
            rom[30705] = 8'h10 ;
            rom[30706] = 8'he6 ;
            rom[30707] = 8'hc6 ;
            rom[30708] = 8'h16 ;
            rom[30709] = 8'hea ;
            rom[30710] = 8'h03 ;
            rom[30711] = 8'h1a ;
            rom[30712] = 8'hdc ;
            rom[30713] = 8'hf0 ;
            rom[30714] = 8'hff ;
            rom[30715] = 8'h2d ;
            rom[30716] = 8'h05 ;
            rom[30717] = 8'h1d ;
            rom[30718] = 8'h0e ;
            rom[30719] = 8'hf9 ;
            rom[30720] = 8'hdc ;
            rom[30721] = 8'hdf ;
            rom[30722] = 8'h03 ;
            rom[30723] = 8'hfd ;
            rom[30724] = 8'hd8 ;
            rom[30725] = 8'hf7 ;
            rom[30726] = 8'h05 ;
            rom[30727] = 8'hfe ;
            rom[30728] = 8'he9 ;
            rom[30729] = 8'he8 ;
            rom[30730] = 8'h1e ;
            rom[30731] = 8'he4 ;
            rom[30732] = 8'hfb ;
            rom[30733] = 8'he3 ;
            rom[30734] = 8'h2c ;
            rom[30735] = 8'hdf ;
            rom[30736] = 8'h0a ;
            rom[30737] = 8'hda ;
            rom[30738] = 8'hea ;
            rom[30739] = 8'h1b ;
            rom[30740] = 8'he1 ;
            rom[30741] = 8'hc4 ;
            rom[30742] = 8'hff ;
            rom[30743] = 8'h06 ;
            rom[30744] = 8'h0e ;
            rom[30745] = 8'he2 ;
            rom[30746] = 8'hff ;
            rom[30747] = 8'hfe ;
            rom[30748] = 8'hf3 ;
            rom[30749] = 8'h08 ;
            rom[30750] = 8'hd2 ;
            rom[30751] = 8'hff ;
            rom[30752] = 8'h01 ;
            rom[30753] = 8'hdf ;
            rom[30754] = 8'h04 ;
            rom[30755] = 8'he1 ;
            rom[30756] = 8'hf1 ;
            rom[30757] = 8'hcf ;
            rom[30758] = 8'he1 ;
            rom[30759] = 8'hf4 ;
            rom[30760] = 8'hef ;
            rom[30761] = 8'h06 ;
            rom[30762] = 8'h19 ;
            rom[30763] = 8'h21 ;
            rom[30764] = 8'h02 ;
            rom[30765] = 8'h0d ;
            rom[30766] = 8'h0a ;
            rom[30767] = 8'hd9 ;
            rom[30768] = 8'hf3 ;
            rom[30769] = 8'hfc ;
            rom[30770] = 8'h06 ;
            rom[30771] = 8'h0b ;
            rom[30772] = 8'hfa ;
            rom[30773] = 8'h0b ;
            rom[30774] = 8'h14 ;
            rom[30775] = 8'h22 ;
            rom[30776] = 8'hd0 ;
            rom[30777] = 8'h0f ;
            rom[30778] = 8'hfd ;
            rom[30779] = 8'h0a ;
            rom[30780] = 8'he9 ;
            rom[30781] = 8'hd2 ;
            rom[30782] = 8'he1 ;
            rom[30783] = 8'hf3 ;
            rom[30784] = 8'hfa ;
            rom[30785] = 8'hf4 ;
            rom[30786] = 8'h0c ;
            rom[30787] = 8'h0f ;
            rom[30788] = 8'hec ;
            rom[30789] = 8'he8 ;
            rom[30790] = 8'h02 ;
            rom[30791] = 8'h24 ;
            rom[30792] = 8'hdf ;
            rom[30793] = 8'hc4 ;
            rom[30794] = 8'h01 ;
            rom[30795] = 8'hec ;
            rom[30796] = 8'hee ;
            rom[30797] = 8'h0a ;
            rom[30798] = 8'he9 ;
            rom[30799] = 8'hed ;
            rom[30800] = 8'h02 ;
            rom[30801] = 8'hd8 ;
            rom[30802] = 8'hf2 ;
            rom[30803] = 8'hf1 ;
            rom[30804] = 8'he7 ;
            rom[30805] = 8'h22 ;
            rom[30806] = 8'hec ;
            rom[30807] = 8'h16 ;
            rom[30808] = 8'h05 ;
            rom[30809] = 8'h1b ;
            rom[30810] = 8'h1c ;
            rom[30811] = 8'h04 ;
            rom[30812] = 8'hf3 ;
            rom[30813] = 8'hd1 ;
            rom[30814] = 8'h10 ;
            rom[30815] = 8'hfb ;
            rom[30816] = 8'hf4 ;
            rom[30817] = 8'hf0 ;
            rom[30818] = 8'hf5 ;
            rom[30819] = 8'hf2 ;
            rom[30820] = 8'hce ;
            rom[30821] = 8'hfe ;
            rom[30822] = 8'h0a ;
            rom[30823] = 8'h11 ;
            rom[30824] = 8'h17 ;
            rom[30825] = 8'hda ;
            rom[30826] = 8'heb ;
            rom[30827] = 8'h14 ;
            rom[30828] = 8'h09 ;
            rom[30829] = 8'h12 ;
            rom[30830] = 8'he1 ;
            rom[30831] = 8'h18 ;
            rom[30832] = 8'h1e ;
            rom[30833] = 8'h20 ;
            rom[30834] = 8'h0b ;
            rom[30835] = 8'he6 ;
            rom[30836] = 8'hef ;
            rom[30837] = 8'hfd ;
            rom[30838] = 8'h12 ;
            rom[30839] = 8'h0b ;
            rom[30840] = 8'h05 ;
            rom[30841] = 8'hff ;
            rom[30842] = 8'h07 ;
            rom[30843] = 8'hf3 ;
            rom[30844] = 8'h06 ;
            rom[30845] = 8'h0f ;
            rom[30846] = 8'h05 ;
            rom[30847] = 8'h04 ;
            rom[30848] = 8'h1a ;
            rom[30849] = 8'hc3 ;
            rom[30850] = 8'hcd ;
            rom[30851] = 8'hef ;
            rom[30852] = 8'hc6 ;
            rom[30853] = 8'h0b ;
            rom[30854] = 8'h02 ;
            rom[30855] = 8'h13 ;
            rom[30856] = 8'hf6 ;
            rom[30857] = 8'hbb ;
            rom[30858] = 8'h2b ;
            rom[30859] = 8'hfd ;
            rom[30860] = 8'h2b ;
            rom[30861] = 8'h02 ;
            rom[30862] = 8'h0f ;
            rom[30863] = 8'h0f ;
            rom[30864] = 8'hf2 ;
            rom[30865] = 8'h11 ;
            rom[30866] = 8'h01 ;
            rom[30867] = 8'h00 ;
            rom[30868] = 8'he7 ;
            rom[30869] = 8'hfa ;
            rom[30870] = 8'he8 ;
            rom[30871] = 8'h0d ;
            rom[30872] = 8'hf7 ;
            rom[30873] = 8'hd4 ;
            rom[30874] = 8'h0a ;
            rom[30875] = 8'hfe ;
            rom[30876] = 8'hf5 ;
            rom[30877] = 8'hf6 ;
            rom[30878] = 8'hf1 ;
            rom[30879] = 8'h03 ;
            rom[30880] = 8'hee ;
            rom[30881] = 8'h01 ;
            rom[30882] = 8'h14 ;
            rom[30883] = 8'hfe ;
            rom[30884] = 8'hf7 ;
            rom[30885] = 8'he9 ;
            rom[30886] = 8'h06 ;
            rom[30887] = 8'hdd ;
            rom[30888] = 8'hf7 ;
            rom[30889] = 8'he5 ;
            rom[30890] = 8'h1c ;
            rom[30891] = 8'h15 ;
            rom[30892] = 8'hf0 ;
            rom[30893] = 8'h09 ;
            rom[30894] = 8'h1e ;
            rom[30895] = 8'hd9 ;
            rom[30896] = 8'he9 ;
            rom[30897] = 8'hdf ;
            rom[30898] = 8'hf6 ;
            rom[30899] = 8'h0d ;
            rom[30900] = 8'hf5 ;
            rom[30901] = 8'h05 ;
            rom[30902] = 8'hff ;
            rom[30903] = 8'h13 ;
            rom[30904] = 8'he7 ;
            rom[30905] = 8'h00 ;
            rom[30906] = 8'h01 ;
            rom[30907] = 8'hed ;
            rom[30908] = 8'hed ;
            rom[30909] = 8'hfb ;
            rom[30910] = 8'h05 ;
            rom[30911] = 8'h24 ;
            rom[30912] = 8'hdf ;
            rom[30913] = 8'h03 ;
            rom[30914] = 8'hee ;
            rom[30915] = 8'hdd ;
            rom[30916] = 8'hff ;
            rom[30917] = 8'h1f ;
            rom[30918] = 8'h03 ;
            rom[30919] = 8'hec ;
            rom[30920] = 8'hed ;
            rom[30921] = 8'hcf ;
            rom[30922] = 8'hd6 ;
            rom[30923] = 8'hde ;
            rom[30924] = 8'hcd ;
            rom[30925] = 8'h01 ;
            rom[30926] = 8'hf6 ;
            rom[30927] = 8'h09 ;
            rom[30928] = 8'h01 ;
            rom[30929] = 8'hf1 ;
            rom[30930] = 8'h08 ;
            rom[30931] = 8'he6 ;
            rom[30932] = 8'h0e ;
            rom[30933] = 8'hf3 ;
            rom[30934] = 8'hd6 ;
            rom[30935] = 8'h1b ;
            rom[30936] = 8'hd4 ;
            rom[30937] = 8'hec ;
            rom[30938] = 8'h1d ;
            rom[30939] = 8'h05 ;
            rom[30940] = 8'h0a ;
            rom[30941] = 8'hf2 ;
            rom[30942] = 8'h0f ;
            rom[30943] = 8'hef ;
            rom[30944] = 8'hc2 ;
            rom[30945] = 8'h0e ;
            rom[30946] = 8'hd1 ;
            rom[30947] = 8'heb ;
            rom[30948] = 8'hc0 ;
            rom[30949] = 8'hd6 ;
            rom[30950] = 8'hf1 ;
            rom[30951] = 8'hfa ;
            rom[30952] = 8'h0a ;
            rom[30953] = 8'hf0 ;
            rom[30954] = 8'h14 ;
            rom[30955] = 8'h0b ;
            rom[30956] = 8'hed ;
            rom[30957] = 8'he8 ;
            rom[30958] = 8'hf8 ;
            rom[30959] = 8'h00 ;
            rom[30960] = 8'h01 ;
            rom[30961] = 8'h25 ;
            rom[30962] = 8'hf4 ;
            rom[30963] = 8'hf3 ;
            rom[30964] = 8'h0d ;
            rom[30965] = 8'hfb ;
            rom[30966] = 8'hfa ;
            rom[30967] = 8'h00 ;
            rom[30968] = 8'h12 ;
            rom[30969] = 8'hf4 ;
            rom[30970] = 8'hd9 ;
            rom[30971] = 8'hed ;
            rom[30972] = 8'hd3 ;
            rom[30973] = 8'h0b ;
            rom[30974] = 8'he6 ;
            rom[30975] = 8'hd3 ;
            rom[30976] = 8'h08 ;
            rom[30977] = 8'h0b ;
            rom[30978] = 8'h04 ;
            rom[30979] = 8'hd0 ;
            rom[30980] = 8'hf6 ;
            rom[30981] = 8'hea ;
            rom[30982] = 8'h20 ;
            rom[30983] = 8'h02 ;
            rom[30984] = 8'hf0 ;
            rom[30985] = 8'h0e ;
            rom[30986] = 8'hcb ;
            rom[30987] = 8'h0a ;
            rom[30988] = 8'h15 ;
            rom[30989] = 8'h12 ;
            rom[30990] = 8'hd9 ;
            rom[30991] = 8'h0a ;
            rom[30992] = 8'hf3 ;
            rom[30993] = 8'h09 ;
            rom[30994] = 8'hdf ;
            rom[30995] = 8'hf2 ;
            rom[30996] = 8'he1 ;
            rom[30997] = 8'h2a ;
            rom[30998] = 8'h07 ;
            rom[30999] = 8'hf7 ;
            rom[31000] = 8'hc7 ;
            rom[31001] = 8'h08 ;
            rom[31002] = 8'hfd ;
            rom[31003] = 8'h05 ;
            rom[31004] = 8'he5 ;
            rom[31005] = 8'hf8 ;
            rom[31006] = 8'hd1 ;
            rom[31007] = 8'hf3 ;
            rom[31008] = 8'h03 ;
            rom[31009] = 8'h13 ;
            rom[31010] = 8'hf3 ;
            rom[31011] = 8'h14 ;
            rom[31012] = 8'h17 ;
            rom[31013] = 8'he9 ;
            rom[31014] = 8'h17 ;
            rom[31015] = 8'he8 ;
            rom[31016] = 8'h17 ;
            rom[31017] = 8'hdd ;
            rom[31018] = 8'h1c ;
            rom[31019] = 8'hd8 ;
            rom[31020] = 8'h11 ;
            rom[31021] = 8'hec ;
            rom[31022] = 8'h13 ;
            rom[31023] = 8'hcf ;
            rom[31024] = 8'hce ;
            rom[31025] = 8'hef ;
            rom[31026] = 8'h09 ;
            rom[31027] = 8'hf0 ;
            rom[31028] = 8'hfc ;
            rom[31029] = 8'hb8 ;
            rom[31030] = 8'h06 ;
            rom[31031] = 8'hfd ;
            rom[31032] = 8'hf2 ;
            rom[31033] = 8'hfe ;
            rom[31034] = 8'hf6 ;
            rom[31035] = 8'h2c ;
            rom[31036] = 8'h2b ;
            rom[31037] = 8'he7 ;
            rom[31038] = 8'h02 ;
            rom[31039] = 8'hdf ;
            rom[31040] = 8'hf9 ;
            rom[31041] = 8'heb ;
            rom[31042] = 8'hfd ;
            rom[31043] = 8'he3 ;
            rom[31044] = 8'hba ;
            rom[31045] = 8'hfe ;
            rom[31046] = 8'hc8 ;
            rom[31047] = 8'hfb ;
            rom[31048] = 8'hd8 ;
            rom[31049] = 8'h20 ;
            rom[31050] = 8'h10 ;
            rom[31051] = 8'h0a ;
            rom[31052] = 8'hfb ;
            rom[31053] = 8'hfb ;
            rom[31054] = 8'h17 ;
            rom[31055] = 8'h07 ;
            rom[31056] = 8'hb7 ;
            rom[31057] = 8'h0f ;
            rom[31058] = 8'he3 ;
            rom[31059] = 8'hf9 ;
            rom[31060] = 8'h17 ;
            rom[31061] = 8'hf3 ;
            rom[31062] = 8'hee ;
            rom[31063] = 8'hff ;
            rom[31064] = 8'hf5 ;
            rom[31065] = 8'h1e ;
            rom[31066] = 8'h18 ;
            rom[31067] = 8'hf1 ;
            rom[31068] = 8'hfc ;
            rom[31069] = 8'hf6 ;
            rom[31070] = 8'hf6 ;
            rom[31071] = 8'h0e ;
            rom[31072] = 8'hf8 ;
            rom[31073] = 8'hf5 ;
            rom[31074] = 8'hc8 ;
            rom[31075] = 8'h06 ;
            rom[31076] = 8'h36 ;
            rom[31077] = 8'hec ;
            rom[31078] = 8'hea ;
            rom[31079] = 8'h0c ;
            rom[31080] = 8'he8 ;
            rom[31081] = 8'h09 ;
            rom[31082] = 8'he5 ;
            rom[31083] = 8'h18 ;
            rom[31084] = 8'hcb ;
            rom[31085] = 8'h0d ;
            rom[31086] = 8'h0a ;
            rom[31087] = 8'h02 ;
            rom[31088] = 8'hf3 ;
            rom[31089] = 8'h06 ;
            rom[31090] = 8'hff ;
            rom[31091] = 8'h07 ;
            rom[31092] = 8'h08 ;
            rom[31093] = 8'h0c ;
            rom[31094] = 8'h11 ;
            rom[31095] = 8'hf5 ;
            rom[31096] = 8'hfd ;
            rom[31097] = 8'hfa ;
            rom[31098] = 8'hd9 ;
            rom[31099] = 8'h17 ;
            rom[31100] = 8'hf0 ;
            rom[31101] = 8'hdd ;
            rom[31102] = 8'hda ;
            rom[31103] = 8'he9 ;
            rom[31104] = 8'h17 ;
            rom[31105] = 8'h0b ;
            rom[31106] = 8'hff ;
            rom[31107] = 8'h00 ;
            rom[31108] = 8'hfa ;
            rom[31109] = 8'h05 ;
            rom[31110] = 8'hce ;
            rom[31111] = 8'h12 ;
            rom[31112] = 8'h0b ;
            rom[31113] = 8'h21 ;
            rom[31114] = 8'h1e ;
            rom[31115] = 8'hfd ;
            rom[31116] = 8'hee ;
            rom[31117] = 8'hf3 ;
            rom[31118] = 8'h07 ;
            rom[31119] = 8'h17 ;
            rom[31120] = 8'h1e ;
            rom[31121] = 8'hea ;
            rom[31122] = 8'h09 ;
            rom[31123] = 8'he7 ;
            rom[31124] = 8'hea ;
            rom[31125] = 8'he3 ;
            rom[31126] = 8'h24 ;
            rom[31127] = 8'hd7 ;
            rom[31128] = 8'h03 ;
            rom[31129] = 8'h03 ;
            rom[31130] = 8'hdb ;
            rom[31131] = 8'hff ;
            rom[31132] = 8'h0e ;
            rom[31133] = 8'h17 ;
            rom[31134] = 8'hd9 ;
            rom[31135] = 8'hdd ;
            rom[31136] = 8'h19 ;
            rom[31137] = 8'h0a ;
            rom[31138] = 8'hff ;
            rom[31139] = 8'h22 ;
            rom[31140] = 8'he8 ;
            rom[31141] = 8'h08 ;
            rom[31142] = 8'hea ;
            rom[31143] = 8'h00 ;
            rom[31144] = 8'h19 ;
            rom[31145] = 8'hf6 ;
            rom[31146] = 8'h04 ;
            rom[31147] = 8'h08 ;
            rom[31148] = 8'hdf ;
            rom[31149] = 8'he4 ;
            rom[31150] = 8'hf7 ;
            rom[31151] = 8'hfe ;
            rom[31152] = 8'hf3 ;
            rom[31153] = 8'he5 ;
            rom[31154] = 8'h23 ;
            rom[31155] = 8'h08 ;
            rom[31156] = 8'he1 ;
            rom[31157] = 8'h15 ;
            rom[31158] = 8'h15 ;
            rom[31159] = 8'had ;
            rom[31160] = 8'hfc ;
            rom[31161] = 8'hfc ;
            rom[31162] = 8'h19 ;
            rom[31163] = 8'he8 ;
            rom[31164] = 8'h23 ;
            rom[31165] = 8'hd1 ;
            rom[31166] = 8'h17 ;
            rom[31167] = 8'h14 ;
            rom[31168] = 8'hdf ;
            rom[31169] = 8'h14 ;
            rom[31170] = 8'h0a ;
            rom[31171] = 8'h01 ;
            rom[31172] = 8'hc2 ;
            rom[31173] = 8'hfb ;
            rom[31174] = 8'hf6 ;
            rom[31175] = 8'h07 ;
            rom[31176] = 8'h06 ;
            rom[31177] = 8'hd4 ;
            rom[31178] = 8'he1 ;
            rom[31179] = 8'he3 ;
            rom[31180] = 8'hf0 ;
            rom[31181] = 8'he8 ;
            rom[31182] = 8'h0a ;
            rom[31183] = 8'hf5 ;
            rom[31184] = 8'h1e ;
            rom[31185] = 8'he7 ;
            rom[31186] = 8'h15 ;
            rom[31187] = 8'he3 ;
            rom[31188] = 8'h16 ;
            rom[31189] = 8'hee ;
            rom[31190] = 8'he1 ;
            rom[31191] = 8'he0 ;
            rom[31192] = 8'h0d ;
            rom[31193] = 8'heb ;
            rom[31194] = 8'h27 ;
            rom[31195] = 8'hff ;
            rom[31196] = 8'hfb ;
            rom[31197] = 8'hdd ;
            rom[31198] = 8'h0c ;
            rom[31199] = 8'h10 ;
            rom[31200] = 8'he7 ;
            rom[31201] = 8'h14 ;
            rom[31202] = 8'hf5 ;
            rom[31203] = 8'he8 ;
            rom[31204] = 8'hf2 ;
            rom[31205] = 8'hd0 ;
            rom[31206] = 8'h04 ;
            rom[31207] = 8'h06 ;
            rom[31208] = 8'hd8 ;
            rom[31209] = 8'h1f ;
            rom[31210] = 8'hea ;
            rom[31211] = 8'h0c ;
            rom[31212] = 8'hf7 ;
            rom[31213] = 8'h15 ;
            rom[31214] = 8'he4 ;
            rom[31215] = 8'hdf ;
            rom[31216] = 8'h05 ;
            rom[31217] = 8'h09 ;
            rom[31218] = 8'hf3 ;
            rom[31219] = 8'h0e ;
            rom[31220] = 8'h07 ;
            rom[31221] = 8'hff ;
            rom[31222] = 8'h04 ;
            rom[31223] = 8'h20 ;
            rom[31224] = 8'h07 ;
            rom[31225] = 8'h02 ;
            rom[31226] = 8'h0e ;
            rom[31227] = 8'hc5 ;
            rom[31228] = 8'he9 ;
            rom[31229] = 8'hec ;
            rom[31230] = 8'hf8 ;
            rom[31231] = 8'hf7 ;
            rom[31232] = 8'h02 ;
            rom[31233] = 8'hf5 ;
            rom[31234] = 8'hd5 ;
            rom[31235] = 8'h08 ;
            rom[31236] = 8'h28 ;
            rom[31237] = 8'h04 ;
            rom[31238] = 8'he8 ;
            rom[31239] = 8'h25 ;
            rom[31240] = 8'h05 ;
            rom[31241] = 8'h06 ;
            rom[31242] = 8'h01 ;
            rom[31243] = 8'h02 ;
            rom[31244] = 8'hd7 ;
            rom[31245] = 8'he5 ;
            rom[31246] = 8'hf4 ;
            rom[31247] = 8'hf9 ;
            rom[31248] = 8'h04 ;
            rom[31249] = 8'hd4 ;
            rom[31250] = 8'h35 ;
            rom[31251] = 8'he4 ;
            rom[31252] = 8'h1f ;
            rom[31253] = 8'he4 ;
            rom[31254] = 8'h10 ;
            rom[31255] = 8'h06 ;
            rom[31256] = 8'hec ;
            rom[31257] = 8'h12 ;
            rom[31258] = 8'h14 ;
            rom[31259] = 8'he6 ;
            rom[31260] = 8'hf2 ;
            rom[31261] = 8'h16 ;
            rom[31262] = 8'hfc ;
            rom[31263] = 8'hba ;
            rom[31264] = 8'h2d ;
            rom[31265] = 8'h03 ;
            rom[31266] = 8'he7 ;
            rom[31267] = 8'h19 ;
            rom[31268] = 8'h01 ;
            rom[31269] = 8'h0f ;
            rom[31270] = 8'h0c ;
            rom[31271] = 8'h0a ;
            rom[31272] = 8'h09 ;
            rom[31273] = 8'hf6 ;
            rom[31274] = 8'h14 ;
            rom[31275] = 8'h02 ;
            rom[31276] = 8'hf2 ;
            rom[31277] = 8'h07 ;
            rom[31278] = 8'he9 ;
            rom[31279] = 8'hee ;
            rom[31280] = 8'he5 ;
            rom[31281] = 8'h00 ;
            rom[31282] = 8'h09 ;
            rom[31283] = 8'hd8 ;
            rom[31284] = 8'hdf ;
            rom[31285] = 8'h00 ;
            rom[31286] = 8'h25 ;
            rom[31287] = 8'h05 ;
            rom[31288] = 8'h0b ;
            rom[31289] = 8'h40 ;
            rom[31290] = 8'h0a ;
            rom[31291] = 8'h06 ;
            rom[31292] = 8'hea ;
            rom[31293] = 8'h0d ;
            rom[31294] = 8'hce ;
            rom[31295] = 8'hcd ;
            rom[31296] = 8'h11 ;
            rom[31297] = 8'h04 ;
            rom[31298] = 8'heb ;
            rom[31299] = 8'h10 ;
            rom[31300] = 8'hfd ;
            rom[31301] = 8'hff ;
            rom[31302] = 8'h14 ;
            rom[31303] = 8'hf2 ;
            rom[31304] = 8'he6 ;
            rom[31305] = 8'hf3 ;
            rom[31306] = 8'h21 ;
            rom[31307] = 8'h09 ;
            rom[31308] = 8'hca ;
            rom[31309] = 8'h11 ;
            rom[31310] = 8'hf0 ;
            rom[31311] = 8'h09 ;
            rom[31312] = 8'he4 ;
            rom[31313] = 8'hff ;
            rom[31314] = 8'hec ;
            rom[31315] = 8'hf0 ;
            rom[31316] = 8'hfa ;
            rom[31317] = 8'hdc ;
            rom[31318] = 8'hf1 ;
            rom[31319] = 8'hf2 ;
            rom[31320] = 8'he2 ;
            rom[31321] = 8'h0d ;
            rom[31322] = 8'hef ;
            rom[31323] = 8'hef ;
            rom[31324] = 8'hf6 ;
            rom[31325] = 8'he3 ;
            rom[31326] = 8'hf7 ;
            rom[31327] = 8'h00 ;
            rom[31328] = 8'h1c ;
            rom[31329] = 8'h20 ;
            rom[31330] = 8'h00 ;
            rom[31331] = 8'h1e ;
            rom[31332] = 8'h14 ;
            rom[31333] = 8'h14 ;
            rom[31334] = 8'he3 ;
            rom[31335] = 8'hb9 ;
            rom[31336] = 8'hf1 ;
            rom[31337] = 8'hfa ;
            rom[31338] = 8'hd6 ;
            rom[31339] = 8'h26 ;
            rom[31340] = 8'hf8 ;
            rom[31341] = 8'hed ;
            rom[31342] = 8'h02 ;
            rom[31343] = 8'hfd ;
            rom[31344] = 8'hea ;
            rom[31345] = 8'hb8 ;
            rom[31346] = 8'h19 ;
            rom[31347] = 8'h0a ;
            rom[31348] = 8'he9 ;
            rom[31349] = 8'hf2 ;
            rom[31350] = 8'hcd ;
            rom[31351] = 8'hdc ;
            rom[31352] = 8'h17 ;
            rom[31353] = 8'hfe ;
            rom[31354] = 8'h05 ;
            rom[31355] = 8'hfb ;
            rom[31356] = 8'he6 ;
            rom[31357] = 8'heb ;
            rom[31358] = 8'hd9 ;
            rom[31359] = 8'h22 ;
            rom[31360] = 8'hde ;
            rom[31361] = 8'hff ;
            rom[31362] = 8'heb ;
            rom[31363] = 8'h10 ;
            rom[31364] = 8'hed ;
            rom[31365] = 8'he1 ;
            rom[31366] = 8'h38 ;
            rom[31367] = 8'hfa ;
            rom[31368] = 8'h08 ;
            rom[31369] = 8'hda ;
            rom[31370] = 8'he2 ;
            rom[31371] = 8'hf8 ;
            rom[31372] = 8'he5 ;
            rom[31373] = 8'hf1 ;
            rom[31374] = 8'h13 ;
            rom[31375] = 8'h17 ;
            rom[31376] = 8'he3 ;
            rom[31377] = 8'he6 ;
            rom[31378] = 8'h01 ;
            rom[31379] = 8'h0a ;
            rom[31380] = 8'h1f ;
            rom[31381] = 8'hf4 ;
            rom[31382] = 8'h0b ;
            rom[31383] = 8'h01 ;
            rom[31384] = 8'h1d ;
            rom[31385] = 8'hd8 ;
            rom[31386] = 8'hff ;
            rom[31387] = 8'h12 ;
            rom[31388] = 8'hf5 ;
            rom[31389] = 8'h00 ;
            rom[31390] = 8'h0a ;
            rom[31391] = 8'hf9 ;
            rom[31392] = 8'h05 ;
            rom[31393] = 8'h11 ;
            rom[31394] = 8'h0f ;
            rom[31395] = 8'hc8 ;
            rom[31396] = 8'hf8 ;
            rom[31397] = 8'heb ;
            rom[31398] = 8'he5 ;
            rom[31399] = 8'h13 ;
            rom[31400] = 8'h04 ;
            rom[31401] = 8'h02 ;
            rom[31402] = 8'h16 ;
            rom[31403] = 8'h13 ;
            rom[31404] = 8'h0b ;
            rom[31405] = 8'hf0 ;
            rom[31406] = 8'hf2 ;
            rom[31407] = 8'hf7 ;
            rom[31408] = 8'hff ;
            rom[31409] = 8'h1d ;
            rom[31410] = 8'h03 ;
            rom[31411] = 8'hef ;
            rom[31412] = 8'hfc ;
            rom[31413] = 8'h04 ;
            rom[31414] = 8'he0 ;
            rom[31415] = 8'h12 ;
            rom[31416] = 8'h0b ;
            rom[31417] = 8'hd9 ;
            rom[31418] = 8'h00 ;
            rom[31419] = 8'h13 ;
            rom[31420] = 8'hf7 ;
            rom[31421] = 8'h18 ;
            rom[31422] = 8'h05 ;
            rom[31423] = 8'hca ;
            rom[31424] = 8'h29 ;
            rom[31425] = 8'h10 ;
            rom[31426] = 8'heb ;
            rom[31427] = 8'hd6 ;
            rom[31428] = 8'h08 ;
            rom[31429] = 8'h08 ;
            rom[31430] = 8'hee ;
            rom[31431] = 8'hd8 ;
            rom[31432] = 8'h18 ;
            rom[31433] = 8'he8 ;
            rom[31434] = 8'hf8 ;
            rom[31435] = 8'h1d ;
            rom[31436] = 8'he5 ;
            rom[31437] = 8'h1c ;
            rom[31438] = 8'heb ;
            rom[31439] = 8'h16 ;
            rom[31440] = 8'h09 ;
            rom[31441] = 8'h10 ;
            rom[31442] = 8'hfd ;
            rom[31443] = 8'hf2 ;
            rom[31444] = 8'hf9 ;
            rom[31445] = 8'heb ;
            rom[31446] = 8'h04 ;
            rom[31447] = 8'he2 ;
            rom[31448] = 8'h16 ;
            rom[31449] = 8'h1c ;
            rom[31450] = 8'hfb ;
            rom[31451] = 8'hdd ;
            rom[31452] = 8'h15 ;
            rom[31453] = 8'h1e ;
            rom[31454] = 8'he7 ;
            rom[31455] = 8'he3 ;
            rom[31456] = 8'hfa ;
            rom[31457] = 8'h18 ;
            rom[31458] = 8'hf9 ;
            rom[31459] = 8'h12 ;
            rom[31460] = 8'hea ;
            rom[31461] = 8'h1f ;
            rom[31462] = 8'h04 ;
            rom[31463] = 8'he2 ;
            rom[31464] = 8'h0c ;
            rom[31465] = 8'hd1 ;
            rom[31466] = 8'hf7 ;
            rom[31467] = 8'h07 ;
            rom[31468] = 8'hd7 ;
            rom[31469] = 8'he1 ;
            rom[31470] = 8'he1 ;
            rom[31471] = 8'h1d ;
            rom[31472] = 8'h05 ;
            rom[31473] = 8'h20 ;
            rom[31474] = 8'he4 ;
            rom[31475] = 8'he6 ;
            rom[31476] = 8'h1c ;
            rom[31477] = 8'h0b ;
            rom[31478] = 8'h11 ;
            rom[31479] = 8'hfe ;
            rom[31480] = 8'hf9 ;
            rom[31481] = 8'h03 ;
            rom[31482] = 8'hc7 ;
            rom[31483] = 8'h25 ;
            rom[31484] = 8'he9 ;
            rom[31485] = 8'h26 ;
            rom[31486] = 8'hc9 ;
            rom[31487] = 8'hfa ;
            rom[31488] = 8'he0 ;
            rom[31489] = 8'hce ;
            rom[31490] = 8'h1c ;
            rom[31491] = 8'heb ;
            rom[31492] = 8'h10 ;
            rom[31493] = 8'h14 ;
            rom[31494] = 8'hc2 ;
            rom[31495] = 8'h09 ;
            rom[31496] = 8'h03 ;
            rom[31497] = 8'hef ;
            rom[31498] = 8'h02 ;
            rom[31499] = 8'h02 ;
            rom[31500] = 8'he3 ;
            rom[31501] = 8'h25 ;
            rom[31502] = 8'h04 ;
            rom[31503] = 8'hfd ;
            rom[31504] = 8'hfa ;
            rom[31505] = 8'h02 ;
            rom[31506] = 8'hd8 ;
            rom[31507] = 8'he3 ;
            rom[31508] = 8'he5 ;
            rom[31509] = 8'h0c ;
            rom[31510] = 8'h2b ;
            rom[31511] = 8'hc2 ;
            rom[31512] = 8'hf1 ;
            rom[31513] = 8'h11 ;
            rom[31514] = 8'hfb ;
            rom[31515] = 8'h37 ;
            rom[31516] = 8'h26 ;
            rom[31517] = 8'hff ;
            rom[31518] = 8'he4 ;
            rom[31519] = 8'hde ;
            rom[31520] = 8'hf8 ;
            rom[31521] = 8'hf8 ;
            rom[31522] = 8'he6 ;
            rom[31523] = 8'h19 ;
            rom[31524] = 8'h11 ;
            rom[31525] = 8'hb6 ;
            rom[31526] = 8'hf4 ;
            rom[31527] = 8'hd6 ;
            rom[31528] = 8'h01 ;
            rom[31529] = 8'hff ;
            rom[31530] = 8'h12 ;
            rom[31531] = 8'hd8 ;
            rom[31532] = 8'hde ;
            rom[31533] = 8'hf7 ;
            rom[31534] = 8'hee ;
            rom[31535] = 8'h15 ;
            rom[31536] = 8'hfa ;
            rom[31537] = 8'hf0 ;
            rom[31538] = 8'h12 ;
            rom[31539] = 8'hdc ;
            rom[31540] = 8'he5 ;
            rom[31541] = 8'h0f ;
            rom[31542] = 8'h09 ;
            rom[31543] = 8'h00 ;
            rom[31544] = 8'hf9 ;
            rom[31545] = 8'h2c ;
            rom[31546] = 8'hf8 ;
            rom[31547] = 8'hf7 ;
            rom[31548] = 8'h02 ;
            rom[31549] = 8'hee ;
            rom[31550] = 8'he1 ;
            rom[31551] = 8'h0a ;
            rom[31552] = 8'h13 ;
            rom[31553] = 8'h03 ;
            rom[31554] = 8'hf9 ;
            rom[31555] = 8'he9 ;
            rom[31556] = 8'hfe ;
            rom[31557] = 8'he6 ;
            rom[31558] = 8'h1f ;
            rom[31559] = 8'h14 ;
            rom[31560] = 8'h08 ;
            rom[31561] = 8'he0 ;
            rom[31562] = 8'h19 ;
            rom[31563] = 8'h10 ;
            rom[31564] = 8'h1c ;
            rom[31565] = 8'h17 ;
            rom[31566] = 8'h0f ;
            rom[31567] = 8'h26 ;
            rom[31568] = 8'h12 ;
            rom[31569] = 8'h0c ;
            rom[31570] = 8'he8 ;
            rom[31571] = 8'hfe ;
            rom[31572] = 8'hf0 ;
            rom[31573] = 8'hf8 ;
            rom[31574] = 8'h10 ;
            rom[31575] = 8'h22 ;
            rom[31576] = 8'h05 ;
            rom[31577] = 8'h06 ;
            rom[31578] = 8'hfc ;
            rom[31579] = 8'h0c ;
            rom[31580] = 8'h06 ;
            rom[31581] = 8'he6 ;
            rom[31582] = 8'h02 ;
            rom[31583] = 8'hf1 ;
            rom[31584] = 8'he1 ;
            rom[31585] = 8'hf6 ;
            rom[31586] = 8'hde ;
            rom[31587] = 8'hcd ;
            rom[31588] = 8'hec ;
            rom[31589] = 8'hee ;
            rom[31590] = 8'hf4 ;
            rom[31591] = 8'h28 ;
            rom[31592] = 8'hdd ;
            rom[31593] = 8'h0e ;
            rom[31594] = 8'h0a ;
            rom[31595] = 8'h05 ;
            rom[31596] = 8'hf4 ;
            rom[31597] = 8'hf9 ;
            rom[31598] = 8'hfd ;
            rom[31599] = 8'h0b ;
            rom[31600] = 8'hf5 ;
            rom[31601] = 8'h25 ;
            rom[31602] = 8'h21 ;
            rom[31603] = 8'hef ;
            rom[31604] = 8'hf7 ;
            rom[31605] = 8'hf5 ;
            rom[31606] = 8'h17 ;
            rom[31607] = 8'h06 ;
            rom[31608] = 8'h18 ;
            rom[31609] = 8'hf7 ;
            rom[31610] = 8'h07 ;
            rom[31611] = 8'hf7 ;
            rom[31612] = 8'hcf ;
            rom[31613] = 8'hf5 ;
            rom[31614] = 8'h1f ;
            rom[31615] = 8'h9d ;
            rom[31616] = 8'hf8 ;
            rom[31617] = 8'h0c ;
            rom[31618] = 8'h00 ;
            rom[31619] = 8'h06 ;
            rom[31620] = 8'h05 ;
            rom[31621] = 8'hcb ;
            rom[31622] = 8'hf3 ;
            rom[31623] = 8'he8 ;
            rom[31624] = 8'hfa ;
            rom[31625] = 8'hf8 ;
            rom[31626] = 8'h09 ;
            rom[31627] = 8'h0a ;
            rom[31628] = 8'hd2 ;
            rom[31629] = 8'hf3 ;
            rom[31630] = 8'hea ;
            rom[31631] = 8'h00 ;
            rom[31632] = 8'hde ;
            rom[31633] = 8'h0a ;
            rom[31634] = 8'h0d ;
            rom[31635] = 8'he2 ;
            rom[31636] = 8'hf4 ;
            rom[31637] = 8'hfe ;
            rom[31638] = 8'hcc ;
            rom[31639] = 8'hfe ;
            rom[31640] = 8'h00 ;
            rom[31641] = 8'h07 ;
            rom[31642] = 8'h26 ;
            rom[31643] = 8'h17 ;
            rom[31644] = 8'hb3 ;
            rom[31645] = 8'hf0 ;
            rom[31646] = 8'h02 ;
            rom[31647] = 8'h0c ;
            rom[31648] = 8'h12 ;
            rom[31649] = 8'hee ;
            rom[31650] = 8'hee ;
            rom[31651] = 8'h01 ;
            rom[31652] = 8'hfa ;
            rom[31653] = 8'hfc ;
            rom[31654] = 8'h1c ;
            rom[31655] = 8'h13 ;
            rom[31656] = 8'h0d ;
            rom[31657] = 8'hfc ;
            rom[31658] = 8'h01 ;
            rom[31659] = 8'he8 ;
            rom[31660] = 8'hda ;
            rom[31661] = 8'h09 ;
            rom[31662] = 8'hff ;
            rom[31663] = 8'he3 ;
            rom[31664] = 8'he2 ;
            rom[31665] = 8'h17 ;
            rom[31666] = 8'h2b ;
            rom[31667] = 8'hcd ;
            rom[31668] = 8'hf5 ;
            rom[31669] = 8'he4 ;
            rom[31670] = 8'hfa ;
            rom[31671] = 8'h1d ;
            rom[31672] = 8'h20 ;
            rom[31673] = 8'he9 ;
            rom[31674] = 8'h20 ;
            rom[31675] = 8'h02 ;
            rom[31676] = 8'h01 ;
            rom[31677] = 8'hf4 ;
            rom[31678] = 8'h16 ;
            rom[31679] = 8'hc6 ;
            rom[31680] = 8'h22 ;
            rom[31681] = 8'he0 ;
            rom[31682] = 8'hf1 ;
            rom[31683] = 8'heb ;
            rom[31684] = 8'hf6 ;
            rom[31685] = 8'h2c ;
            rom[31686] = 8'hd5 ;
            rom[31687] = 8'he1 ;
            rom[31688] = 8'hfb ;
            rom[31689] = 8'h05 ;
            rom[31690] = 8'hf5 ;
            rom[31691] = 8'hda ;
            rom[31692] = 8'h11 ;
            rom[31693] = 8'hf0 ;
            rom[31694] = 8'h06 ;
            rom[31695] = 8'h07 ;
            rom[31696] = 8'hb7 ;
            rom[31697] = 8'h0c ;
            rom[31698] = 8'hea ;
            rom[31699] = 8'hfb ;
            rom[31700] = 8'hee ;
            rom[31701] = 8'hd5 ;
            rom[31702] = 8'h0d ;
            rom[31703] = 8'h0d ;
            rom[31704] = 8'heb ;
            rom[31705] = 8'h19 ;
            rom[31706] = 8'he7 ;
            rom[31707] = 8'hdc ;
            rom[31708] = 8'hfb ;
            rom[31709] = 8'h1f ;
            rom[31710] = 8'h14 ;
            rom[31711] = 8'hf4 ;
            rom[31712] = 8'hf6 ;
            rom[31713] = 8'hdc ;
            rom[31714] = 8'he2 ;
            rom[31715] = 8'h0d ;
            rom[31716] = 8'h08 ;
            rom[31717] = 8'hf4 ;
            rom[31718] = 8'hf6 ;
            rom[31719] = 8'hb3 ;
            rom[31720] = 8'hfd ;
            rom[31721] = 8'hf8 ;
            rom[31722] = 8'hd3 ;
            rom[31723] = 8'h0f ;
            rom[31724] = 8'hac ;
            rom[31725] = 8'hec ;
            rom[31726] = 8'h01 ;
            rom[31727] = 8'h05 ;
            rom[31728] = 8'hec ;
            rom[31729] = 8'h05 ;
            rom[31730] = 8'h14 ;
            rom[31731] = 8'hf9 ;
            rom[31732] = 8'h04 ;
            rom[31733] = 8'h03 ;
            rom[31734] = 8'h0a ;
            rom[31735] = 8'hd1 ;
            rom[31736] = 8'he1 ;
            rom[31737] = 8'he3 ;
            rom[31738] = 8'he1 ;
            rom[31739] = 8'h12 ;
            rom[31740] = 8'hfd ;
            rom[31741] = 8'h05 ;
            rom[31742] = 8'hdc ;
            rom[31743] = 8'hd6 ;
            rom[31744] = 8'hf4 ;
            rom[31745] = 8'hf5 ;
            rom[31746] = 8'hec ;
            rom[31747] = 8'hed ;
            rom[31748] = 8'h04 ;
            rom[31749] = 8'hff ;
            rom[31750] = 8'h15 ;
            rom[31751] = 8'h03 ;
            rom[31752] = 8'h11 ;
            rom[31753] = 8'hda ;
            rom[31754] = 8'h03 ;
            rom[31755] = 8'hf5 ;
            rom[31756] = 8'h0f ;
            rom[31757] = 8'h01 ;
            rom[31758] = 8'hf4 ;
            rom[31759] = 8'h28 ;
            rom[31760] = 8'hec ;
            rom[31761] = 8'he5 ;
            rom[31762] = 8'h24 ;
            rom[31763] = 8'hfc ;
            rom[31764] = 8'h06 ;
            rom[31765] = 8'h22 ;
            rom[31766] = 8'h08 ;
            rom[31767] = 8'h27 ;
            rom[31768] = 8'hfd ;
            rom[31769] = 8'hff ;
            rom[31770] = 8'h0b ;
            rom[31771] = 8'hd9 ;
            rom[31772] = 8'hcb ;
            rom[31773] = 8'h0a ;
            rom[31774] = 8'he4 ;
            rom[31775] = 8'hf8 ;
            rom[31776] = 8'hdc ;
            rom[31777] = 8'h06 ;
            rom[31778] = 8'hfd ;
            rom[31779] = 8'hf0 ;
            rom[31780] = 8'he5 ;
            rom[31781] = 8'hf6 ;
            rom[31782] = 8'h0b ;
            rom[31783] = 8'hf9 ;
            rom[31784] = 8'he6 ;
            rom[31785] = 8'hf9 ;
            rom[31786] = 8'hed ;
            rom[31787] = 8'h11 ;
            rom[31788] = 8'he7 ;
            rom[31789] = 8'h1a ;
            rom[31790] = 8'hd5 ;
            rom[31791] = 8'h0e ;
            rom[31792] = 8'hff ;
            rom[31793] = 8'h15 ;
            rom[31794] = 8'h0f ;
            rom[31795] = 8'h06 ;
            rom[31796] = 8'hd0 ;
            rom[31797] = 8'h09 ;
            rom[31798] = 8'h0d ;
            rom[31799] = 8'hf0 ;
            rom[31800] = 8'h0f ;
            rom[31801] = 8'h06 ;
            rom[31802] = 8'h0c ;
            rom[31803] = 8'heb ;
            rom[31804] = 8'h01 ;
            rom[31805] = 8'h07 ;
            rom[31806] = 8'h23 ;
            rom[31807] = 8'hd1 ;
            rom[31808] = 8'hf2 ;
            rom[31809] = 8'h25 ;
            rom[31810] = 8'hdc ;
            rom[31811] = 8'hfa ;
            rom[31812] = 8'he5 ;
            rom[31813] = 8'h1e ;
            rom[31814] = 8'hf6 ;
            rom[31815] = 8'hcf ;
            rom[31816] = 8'h0d ;
            rom[31817] = 8'hfd ;
            rom[31818] = 8'hd0 ;
            rom[31819] = 8'h03 ;
            rom[31820] = 8'hd7 ;
            rom[31821] = 8'h14 ;
            rom[31822] = 8'hda ;
            rom[31823] = 8'hed ;
            rom[31824] = 8'hef ;
            rom[31825] = 8'h2f ;
            rom[31826] = 8'h0c ;
            rom[31827] = 8'hef ;
            rom[31828] = 8'hfd ;
            rom[31829] = 8'hea ;
            rom[31830] = 8'hff ;
            rom[31831] = 8'hf7 ;
            rom[31832] = 8'hef ;
            rom[31833] = 8'h0a ;
            rom[31834] = 8'hf4 ;
            rom[31835] = 8'he7 ;
            rom[31836] = 8'hcc ;
            rom[31837] = 8'hfd ;
            rom[31838] = 8'hf1 ;
            rom[31839] = 8'hca ;
            rom[31840] = 8'hff ;
            rom[31841] = 8'h24 ;
            rom[31842] = 8'hf4 ;
            rom[31843] = 8'h13 ;
            rom[31844] = 8'h07 ;
            rom[31845] = 8'he9 ;
            rom[31846] = 8'hf7 ;
            rom[31847] = 8'hbb ;
            rom[31848] = 8'hfe ;
            rom[31849] = 8'hf6 ;
            rom[31850] = 8'he4 ;
            rom[31851] = 8'h24 ;
            rom[31852] = 8'hf4 ;
            rom[31853] = 8'he8 ;
            rom[31854] = 8'hed ;
            rom[31855] = 8'hd8 ;
            rom[31856] = 8'h02 ;
            rom[31857] = 8'h08 ;
            rom[31858] = 8'hd8 ;
            rom[31859] = 8'hdb ;
            rom[31860] = 8'hfe ;
            rom[31861] = 8'hfe ;
            rom[31862] = 8'hd0 ;
            rom[31863] = 8'hd6 ;
            rom[31864] = 8'h0d ;
            rom[31865] = 8'he6 ;
            rom[31866] = 8'hfa ;
            rom[31867] = 8'h05 ;
            rom[31868] = 8'h1c ;
            rom[31869] = 8'hf4 ;
            rom[31870] = 8'he0 ;
            rom[31871] = 8'hf9 ;
            rom[31872] = 8'hf9 ;
            rom[31873] = 8'hf5 ;
            rom[31874] = 8'hfd ;
            rom[31875] = 8'hf8 ;
            rom[31876] = 8'h09 ;
            rom[31877] = 8'h11 ;
            rom[31878] = 8'hf8 ;
            rom[31879] = 8'h00 ;
            rom[31880] = 8'hec ;
            rom[31881] = 8'h13 ;
            rom[31882] = 8'h1b ;
            rom[31883] = 8'hff ;
            rom[31884] = 8'h0a ;
            rom[31885] = 8'h08 ;
            rom[31886] = 8'hff ;
            rom[31887] = 8'h0b ;
            rom[31888] = 8'hff ;
            rom[31889] = 8'h0e ;
            rom[31890] = 8'hd3 ;
            rom[31891] = 8'he8 ;
            rom[31892] = 8'he3 ;
            rom[31893] = 8'h1b ;
            rom[31894] = 8'h0d ;
            rom[31895] = 8'hd8 ;
            rom[31896] = 8'h01 ;
            rom[31897] = 8'hfc ;
            rom[31898] = 8'h08 ;
            rom[31899] = 8'h19 ;
            rom[31900] = 8'h1b ;
            rom[31901] = 8'he0 ;
            rom[31902] = 8'hcc ;
            rom[31903] = 8'hf8 ;
            rom[31904] = 8'h1b ;
            rom[31905] = 8'h1a ;
            rom[31906] = 8'he2 ;
            rom[31907] = 8'h0e ;
            rom[31908] = 8'hd2 ;
            rom[31909] = 8'hfc ;
            rom[31910] = 8'h02 ;
            rom[31911] = 8'hf6 ;
            rom[31912] = 8'hfe ;
            rom[31913] = 8'h06 ;
            rom[31914] = 8'h14 ;
            rom[31915] = 8'hfd ;
            rom[31916] = 8'h02 ;
            rom[31917] = 8'hd6 ;
            rom[31918] = 8'h00 ;
            rom[31919] = 8'hdf ;
            rom[31920] = 8'hfa ;
            rom[31921] = 8'hfa ;
            rom[31922] = 8'hea ;
            rom[31923] = 8'hfd ;
            rom[31924] = 8'h21 ;
            rom[31925] = 8'hec ;
            rom[31926] = 8'h13 ;
            rom[31927] = 8'he5 ;
            rom[31928] = 8'h01 ;
            rom[31929] = 8'hec ;
            rom[31930] = 8'hee ;
            rom[31931] = 8'h1c ;
            rom[31932] = 8'h01 ;
            rom[31933] = 8'hef ;
            rom[31934] = 8'h01 ;
            rom[31935] = 8'h04 ;
            rom[31936] = 8'h08 ;
            rom[31937] = 8'h04 ;
            rom[31938] = 8'h12 ;
            rom[31939] = 8'hd8 ;
            rom[31940] = 8'he5 ;
            rom[31941] = 8'hf9 ;
            rom[31942] = 8'hee ;
            rom[31943] = 8'h23 ;
            rom[31944] = 8'h04 ;
            rom[31945] = 8'heb ;
            rom[31946] = 8'h07 ;
            rom[31947] = 8'h11 ;
            rom[31948] = 8'h02 ;
            rom[31949] = 8'he9 ;
            rom[31950] = 8'h0b ;
            rom[31951] = 8'h2a ;
            rom[31952] = 8'h14 ;
            rom[31953] = 8'hed ;
            rom[31954] = 8'he7 ;
            rom[31955] = 8'h06 ;
            rom[31956] = 8'he3 ;
            rom[31957] = 8'h06 ;
            rom[31958] = 8'hd5 ;
            rom[31959] = 8'hfd ;
            rom[31960] = 8'h07 ;
            rom[31961] = 8'hea ;
            rom[31962] = 8'h11 ;
            rom[31963] = 8'h0b ;
            rom[31964] = 8'h12 ;
            rom[31965] = 8'hea ;
            rom[31966] = 8'he5 ;
            rom[31967] = 8'h06 ;
            rom[31968] = 8'h02 ;
            rom[31969] = 8'he9 ;
            rom[31970] = 8'h0e ;
            rom[31971] = 8'hef ;
            rom[31972] = 8'h13 ;
            rom[31973] = 8'he4 ;
            rom[31974] = 8'heb ;
            rom[31975] = 8'h1d ;
            rom[31976] = 8'hed ;
            rom[31977] = 8'h09 ;
            rom[31978] = 8'h05 ;
            rom[31979] = 8'h0e ;
            rom[31980] = 8'h02 ;
            rom[31981] = 8'h02 ;
            rom[31982] = 8'hfa ;
            rom[31983] = 8'h26 ;
            rom[31984] = 8'h17 ;
            rom[31985] = 8'h20 ;
            rom[31986] = 8'h05 ;
            rom[31987] = 8'h0e ;
            rom[31988] = 8'h1c ;
            rom[31989] = 8'h07 ;
            rom[31990] = 8'h27 ;
            rom[31991] = 8'h2a ;
            rom[31992] = 8'h0a ;
            rom[31993] = 8'h0e ;
            rom[31994] = 8'h1f ;
            rom[31995] = 8'hdc ;
            rom[31996] = 8'hef ;
            rom[31997] = 8'hf9 ;
            rom[31998] = 8'hf8 ;
            rom[31999] = 8'he8 ;
            rom[32000] = 8'h19 ;
            rom[32001] = 8'hff ;
            rom[32002] = 8'h15 ;
            rom[32003] = 8'he9 ;
            rom[32004] = 8'hf9 ;
            rom[32005] = 8'hed ;
            rom[32006] = 8'he2 ;
            rom[32007] = 8'hfa ;
            rom[32008] = 8'hef ;
            rom[32009] = 8'hfa ;
            rom[32010] = 8'h2b ;
            rom[32011] = 8'ha6 ;
            rom[32012] = 8'hc4 ;
            rom[32013] = 8'hf1 ;
            rom[32014] = 8'h11 ;
            rom[32015] = 8'h15 ;
            rom[32016] = 8'hd0 ;
            rom[32017] = 8'h0f ;
            rom[32018] = 8'he5 ;
            rom[32019] = 8'hdf ;
            rom[32020] = 8'he1 ;
            rom[32021] = 8'hc5 ;
            rom[32022] = 8'h0a ;
            rom[32023] = 8'hed ;
            rom[32024] = 8'hee ;
            rom[32025] = 8'he0 ;
            rom[32026] = 8'hd7 ;
            rom[32027] = 8'hf2 ;
            rom[32028] = 8'h16 ;
            rom[32029] = 8'hf7 ;
            rom[32030] = 8'hf0 ;
            rom[32031] = 8'hf9 ;
            rom[32032] = 8'h01 ;
            rom[32033] = 8'hf9 ;
            rom[32034] = 8'h05 ;
            rom[32035] = 8'h03 ;
            rom[32036] = 8'hef ;
            rom[32037] = 8'hd2 ;
            rom[32038] = 8'he8 ;
            rom[32039] = 8'h20 ;
            rom[32040] = 8'h06 ;
            rom[32041] = 8'h24 ;
            rom[32042] = 8'h09 ;
            rom[32043] = 8'h14 ;
            rom[32044] = 8'hd9 ;
            rom[32045] = 8'hdc ;
            rom[32046] = 8'hee ;
            rom[32047] = 8'hfe ;
            rom[32048] = 8'h0f ;
            rom[32049] = 8'h06 ;
            rom[32050] = 8'hfa ;
            rom[32051] = 8'hed ;
            rom[32052] = 8'hee ;
            rom[32053] = 8'h08 ;
            rom[32054] = 8'h08 ;
            rom[32055] = 8'hea ;
            rom[32056] = 8'h08 ;
            rom[32057] = 8'hec ;
            rom[32058] = 8'hf9 ;
            rom[32059] = 8'hf1 ;
            rom[32060] = 8'hf9 ;
            rom[32061] = 8'hf1 ;
            rom[32062] = 8'hff ;
            rom[32063] = 8'hed ;
            rom[32064] = 8'he1 ;
            rom[32065] = 8'h11 ;
            rom[32066] = 8'hf0 ;
            rom[32067] = 8'hde ;
            rom[32068] = 8'hee ;
            rom[32069] = 8'h1d ;
            rom[32070] = 8'hf8 ;
            rom[32071] = 8'hf7 ;
            rom[32072] = 8'h10 ;
            rom[32073] = 8'h04 ;
            rom[32074] = 8'hf4 ;
            rom[32075] = 8'hd8 ;
            rom[32076] = 8'he4 ;
            rom[32077] = 8'hfa ;
            rom[32078] = 8'h14 ;
            rom[32079] = 8'heb ;
            rom[32080] = 8'h1f ;
            rom[32081] = 8'he8 ;
            rom[32082] = 8'hfd ;
            rom[32083] = 8'hbe ;
            rom[32084] = 8'h02 ;
            rom[32085] = 8'h07 ;
            rom[32086] = 8'hc8 ;
            rom[32087] = 8'h26 ;
            rom[32088] = 8'hf7 ;
            rom[32089] = 8'he4 ;
            rom[32090] = 8'h14 ;
            rom[32091] = 8'h11 ;
            rom[32092] = 8'hfa ;
            rom[32093] = 8'h09 ;
            rom[32094] = 8'hd0 ;
            rom[32095] = 8'hdf ;
            rom[32096] = 8'hd8 ;
            rom[32097] = 8'hea ;
            rom[32098] = 8'h0b ;
            rom[32099] = 8'h00 ;
            rom[32100] = 8'hd9 ;
            rom[32101] = 8'hf8 ;
            rom[32102] = 8'h11 ;
            rom[32103] = 8'h0c ;
            rom[32104] = 8'hcb ;
            rom[32105] = 8'hf8 ;
            rom[32106] = 8'hf8 ;
            rom[32107] = 8'hdb ;
            rom[32108] = 8'h1a ;
            rom[32109] = 8'hfe ;
            rom[32110] = 8'he9 ;
            rom[32111] = 8'h05 ;
            rom[32112] = 8'hea ;
            rom[32113] = 8'h09 ;
            rom[32114] = 8'h08 ;
            rom[32115] = 8'h06 ;
            rom[32116] = 8'hf7 ;
            rom[32117] = 8'h0a ;
            rom[32118] = 8'hf6 ;
            rom[32119] = 8'h0d ;
            rom[32120] = 8'h04 ;
            rom[32121] = 8'heb ;
            rom[32122] = 8'hdd ;
            rom[32123] = 8'hf1 ;
            rom[32124] = 8'hf0 ;
            rom[32125] = 8'hfe ;
            rom[32126] = 8'h1d ;
            rom[32127] = 8'he1 ;
            rom[32128] = 8'h04 ;
            rom[32129] = 8'hf8 ;
            rom[32130] = 8'h04 ;
            rom[32131] = 8'h0c ;
            rom[32132] = 8'h16 ;
            rom[32133] = 8'h06 ;
            rom[32134] = 8'h1a ;
            rom[32135] = 8'h0d ;
            rom[32136] = 8'hf1 ;
            rom[32137] = 8'h09 ;
            rom[32138] = 8'h07 ;
            rom[32139] = 8'hff ;
            rom[32140] = 8'hfe ;
            rom[32141] = 8'hf7 ;
            rom[32142] = 8'h08 ;
            rom[32143] = 8'hfa ;
            rom[32144] = 8'h03 ;
            rom[32145] = 8'hfe ;
            rom[32146] = 8'hef ;
            rom[32147] = 8'hf2 ;
            rom[32148] = 8'h28 ;
            rom[32149] = 8'h11 ;
            rom[32150] = 8'he4 ;
            rom[32151] = 8'hf6 ;
            rom[32152] = 8'hf8 ;
            rom[32153] = 8'h1c ;
            rom[32154] = 8'h11 ;
            rom[32155] = 8'h16 ;
            rom[32156] = 8'hff ;
            rom[32157] = 8'hf0 ;
            rom[32158] = 8'h0f ;
            rom[32159] = 8'h13 ;
            rom[32160] = 8'he4 ;
            rom[32161] = 8'he0 ;
            rom[32162] = 8'hda ;
            rom[32163] = 8'hd5 ;
            rom[32164] = 8'h0c ;
            rom[32165] = 8'hdf ;
            rom[32166] = 8'h09 ;
            rom[32167] = 8'h1b ;
            rom[32168] = 8'h07 ;
            rom[32169] = 8'he7 ;
            rom[32170] = 8'hf4 ;
            rom[32171] = 8'h02 ;
            rom[32172] = 8'h0c ;
            rom[32173] = 8'hd5 ;
            rom[32174] = 8'hfa ;
            rom[32175] = 8'hf6 ;
            rom[32176] = 8'hf3 ;
            rom[32177] = 8'h0b ;
            rom[32178] = 8'h0c ;
            rom[32179] = 8'h08 ;
            rom[32180] = 8'hf8 ;
            rom[32181] = 8'h09 ;
            rom[32182] = 8'hec ;
            rom[32183] = 8'hf4 ;
            rom[32184] = 8'hf5 ;
            rom[32185] = 8'h07 ;
            rom[32186] = 8'h0b ;
            rom[32187] = 8'h0e ;
            rom[32188] = 8'hef ;
            rom[32189] = 8'hfe ;
            rom[32190] = 8'he2 ;
            rom[32191] = 8'hf4 ;
            rom[32192] = 8'h08 ;
            rom[32193] = 8'h0b ;
            rom[32194] = 8'hf9 ;
            rom[32195] = 8'hd7 ;
            rom[32196] = 8'h0d ;
            rom[32197] = 8'he0 ;
            rom[32198] = 8'hfb ;
            rom[32199] = 8'he0 ;
            rom[32200] = 8'h00 ;
            rom[32201] = 8'hf6 ;
            rom[32202] = 8'hfb ;
            rom[32203] = 8'h23 ;
            rom[32204] = 8'h15 ;
            rom[32205] = 8'h0b ;
            rom[32206] = 8'hc5 ;
            rom[32207] = 8'h00 ;
            rom[32208] = 8'hdd ;
            rom[32209] = 8'h0d ;
            rom[32210] = 8'hf8 ;
            rom[32211] = 8'hff ;
            rom[32212] = 8'h14 ;
            rom[32213] = 8'hf9 ;
            rom[32214] = 8'h20 ;
            rom[32215] = 8'h0e ;
            rom[32216] = 8'h08 ;
            rom[32217] = 8'hf1 ;
            rom[32218] = 8'he1 ;
            rom[32219] = 8'h01 ;
            rom[32220] = 8'h0f ;
            rom[32221] = 8'h0e ;
            rom[32222] = 8'hf6 ;
            rom[32223] = 8'he0 ;
            rom[32224] = 8'hea ;
            rom[32225] = 8'he5 ;
            rom[32226] = 8'he4 ;
            rom[32227] = 8'h09 ;
            rom[32228] = 8'h32 ;
            rom[32229] = 8'hcd ;
            rom[32230] = 8'hec ;
            rom[32231] = 8'hdc ;
            rom[32232] = 8'hca ;
            rom[32233] = 8'hdb ;
            rom[32234] = 8'hd9 ;
            rom[32235] = 8'hf5 ;
            rom[32236] = 8'hc1 ;
            rom[32237] = 8'heb ;
            rom[32238] = 8'he1 ;
            rom[32239] = 8'h21 ;
            rom[32240] = 8'h0d ;
            rom[32241] = 8'h09 ;
            rom[32242] = 8'h0d ;
            rom[32243] = 8'hfb ;
            rom[32244] = 8'hf3 ;
            rom[32245] = 8'h06 ;
            rom[32246] = 8'hef ;
            rom[32247] = 8'he8 ;
            rom[32248] = 8'h19 ;
            rom[32249] = 8'hff ;
            rom[32250] = 8'hfd ;
            rom[32251] = 8'h19 ;
            rom[32252] = 8'he5 ;
            rom[32253] = 8'hd7 ;
            rom[32254] = 8'hc2 ;
            rom[32255] = 8'hac ;
            rom[32256] = 8'h0f ;
            rom[32257] = 8'hf5 ;
            rom[32258] = 8'h05 ;
            rom[32259] = 8'hf2 ;
            rom[32260] = 8'hed ;
            rom[32261] = 8'h12 ;
            rom[32262] = 8'hd5 ;
            rom[32263] = 8'h11 ;
            rom[32264] = 8'hcb ;
            rom[32265] = 8'hdf ;
            rom[32266] = 8'h12 ;
            rom[32267] = 8'h02 ;
            rom[32268] = 8'hee ;
            rom[32269] = 8'h0c ;
            rom[32270] = 8'h18 ;
            rom[32271] = 8'hff ;
            rom[32272] = 8'h0a ;
            rom[32273] = 8'h03 ;
            rom[32274] = 8'hcb ;
            rom[32275] = 8'he5 ;
            rom[32276] = 8'hfa ;
            rom[32277] = 8'hea ;
            rom[32278] = 8'hcf ;
            rom[32279] = 8'hf5 ;
            rom[32280] = 8'h17 ;
            rom[32281] = 8'h00 ;
            rom[32282] = 8'h02 ;
            rom[32283] = 8'h0a ;
            rom[32284] = 8'hdc ;
            rom[32285] = 8'hed ;
            rom[32286] = 8'h22 ;
            rom[32287] = 8'hfc ;
            rom[32288] = 8'hff ;
            rom[32289] = 8'h13 ;
            rom[32290] = 8'hdc ;
            rom[32291] = 8'hdc ;
            rom[32292] = 8'h29 ;
            rom[32293] = 8'h05 ;
            rom[32294] = 8'hff ;
            rom[32295] = 8'hf5 ;
            rom[32296] = 8'he0 ;
            rom[32297] = 8'he4 ;
            rom[32298] = 8'hef ;
            rom[32299] = 8'hdf ;
            rom[32300] = 8'h0a ;
            rom[32301] = 8'hd2 ;
            rom[32302] = 8'h04 ;
            rom[32303] = 8'he2 ;
            rom[32304] = 8'hf9 ;
            rom[32305] = 8'hfe ;
            rom[32306] = 8'hf4 ;
            rom[32307] = 8'hce ;
            rom[32308] = 8'h10 ;
            rom[32309] = 8'hd7 ;
            rom[32310] = 8'h17 ;
            rom[32311] = 8'hf5 ;
            rom[32312] = 8'h22 ;
            rom[32313] = 8'hf9 ;
            rom[32314] = 8'h08 ;
            rom[32315] = 8'he3 ;
            rom[32316] = 8'h07 ;
            rom[32317] = 8'he4 ;
            rom[32318] = 8'hed ;
            rom[32319] = 8'h0a ;
            rom[32320] = 8'hf9 ;
            rom[32321] = 8'h0b ;
            rom[32322] = 8'hff ;
            rom[32323] = 8'he2 ;
            rom[32324] = 8'hd3 ;
            rom[32325] = 8'hfd ;
            rom[32326] = 8'hfb ;
            rom[32327] = 8'h0f ;
            rom[32328] = 8'hfd ;
            rom[32329] = 8'h1e ;
            rom[32330] = 8'h05 ;
            rom[32331] = 8'hfa ;
            rom[32332] = 8'hfe ;
            rom[32333] = 8'h21 ;
            rom[32334] = 8'he8 ;
            rom[32335] = 8'h19 ;
            rom[32336] = 8'he8 ;
            rom[32337] = 8'hf5 ;
            rom[32338] = 8'he0 ;
            rom[32339] = 8'h06 ;
            rom[32340] = 8'h0b ;
            rom[32341] = 8'hf1 ;
            rom[32342] = 8'h1e ;
            rom[32343] = 8'h13 ;
            rom[32344] = 8'h0d ;
            rom[32345] = 8'h0c ;
            rom[32346] = 8'hfa ;
            rom[32347] = 8'h13 ;
            rom[32348] = 8'h10 ;
            rom[32349] = 8'hfa ;
            rom[32350] = 8'h1e ;
            rom[32351] = 8'h0d ;
            rom[32352] = 8'h12 ;
            rom[32353] = 8'hd7 ;
            rom[32354] = 8'hef ;
            rom[32355] = 8'hd1 ;
            rom[32356] = 8'hde ;
            rom[32357] = 8'hfe ;
            rom[32358] = 8'h1e ;
            rom[32359] = 8'h00 ;
            rom[32360] = 8'hf2 ;
            rom[32361] = 8'hf1 ;
            rom[32362] = 8'he1 ;
            rom[32363] = 8'he5 ;
            rom[32364] = 8'he2 ;
            rom[32365] = 8'h0a ;
            rom[32366] = 8'h1c ;
            rom[32367] = 8'h1a ;
            rom[32368] = 8'h1d ;
            rom[32369] = 8'h02 ;
            rom[32370] = 8'h08 ;
            rom[32371] = 8'h0f ;
            rom[32372] = 8'h15 ;
            rom[32373] = 8'h11 ;
            rom[32374] = 8'he5 ;
            rom[32375] = 8'h0c ;
            rom[32376] = 8'h01 ;
            rom[32377] = 8'h0d ;
            rom[32378] = 8'h22 ;
            rom[32379] = 8'hfd ;
            rom[32380] = 8'hf0 ;
            rom[32381] = 8'h03 ;
            rom[32382] = 8'hda ;
            rom[32383] = 8'hd7 ;
            rom[32384] = 8'h1d ;
            rom[32385] = 8'h06 ;
            rom[32386] = 8'h03 ;
            rom[32387] = 8'h16 ;
            rom[32388] = 8'h21 ;
            rom[32389] = 8'he7 ;
            rom[32390] = 8'h08 ;
            rom[32391] = 8'h34 ;
            rom[32392] = 8'hfe ;
            rom[32393] = 8'h09 ;
            rom[32394] = 8'h17 ;
            rom[32395] = 8'he3 ;
            rom[32396] = 8'hef ;
            rom[32397] = 8'hd6 ;
            rom[32398] = 8'hf2 ;
            rom[32399] = 8'hfc ;
            rom[32400] = 8'hd2 ;
            rom[32401] = 8'hff ;
            rom[32402] = 8'h21 ;
            rom[32403] = 8'he3 ;
            rom[32404] = 8'h01 ;
            rom[32405] = 8'hd5 ;
            rom[32406] = 8'he2 ;
            rom[32407] = 8'hd6 ;
            rom[32408] = 8'hdb ;
            rom[32409] = 8'h0b ;
            rom[32410] = 8'h05 ;
            rom[32411] = 8'hca ;
            rom[32412] = 8'hfd ;
            rom[32413] = 8'h03 ;
            rom[32414] = 8'h13 ;
            rom[32415] = 8'h08 ;
            rom[32416] = 8'h0e ;
            rom[32417] = 8'h04 ;
            rom[32418] = 8'hef ;
            rom[32419] = 8'h14 ;
            rom[32420] = 8'hcf ;
            rom[32421] = 8'h02 ;
            rom[32422] = 8'hf2 ;
            rom[32423] = 8'h15 ;
            rom[32424] = 8'hfd ;
            rom[32425] = 8'he9 ;
            rom[32426] = 8'he9 ;
            rom[32427] = 8'h08 ;
            rom[32428] = 8'hf9 ;
            rom[32429] = 8'hdf ;
            rom[32430] = 8'hda ;
            rom[32431] = 8'h14 ;
            rom[32432] = 8'hf9 ;
            rom[32433] = 8'hdd ;
            rom[32434] = 8'h01 ;
            rom[32435] = 8'h20 ;
            rom[32436] = 8'hd3 ;
            rom[32437] = 8'h02 ;
            rom[32438] = 8'h10 ;
            rom[32439] = 8'h0c ;
            rom[32440] = 8'h11 ;
            rom[32441] = 8'he8 ;
            rom[32442] = 8'h14 ;
            rom[32443] = 8'hff ;
            rom[32444] = 8'hf7 ;
            rom[32445] = 8'h02 ;
            rom[32446] = 8'h14 ;
            rom[32447] = 8'he2 ;
            rom[32448] = 8'h14 ;
            rom[32449] = 8'h02 ;
            rom[32450] = 8'hf2 ;
            rom[32451] = 8'hcf ;
            rom[32452] = 8'hef ;
            rom[32453] = 8'h0e ;
            rom[32454] = 8'he1 ;
            rom[32455] = 8'he1 ;
            rom[32456] = 8'h0f ;
            rom[32457] = 8'h0b ;
            rom[32458] = 8'hf5 ;
            rom[32459] = 8'h04 ;
            rom[32460] = 8'hf7 ;
            rom[32461] = 8'hed ;
            rom[32462] = 8'hed ;
            rom[32463] = 8'h00 ;
            rom[32464] = 8'h0e ;
            rom[32465] = 8'hf4 ;
            rom[32466] = 8'h1d ;
            rom[32467] = 8'hb5 ;
            rom[32468] = 8'h18 ;
            rom[32469] = 8'hdc ;
            rom[32470] = 8'he5 ;
            rom[32471] = 8'h08 ;
            rom[32472] = 8'h14 ;
            rom[32473] = 8'hf3 ;
            rom[32474] = 8'h19 ;
            rom[32475] = 8'h1a ;
            rom[32476] = 8'h04 ;
            rom[32477] = 8'he0 ;
            rom[32478] = 8'hed ;
            rom[32479] = 8'h0a ;
            rom[32480] = 8'hdd ;
            rom[32481] = 8'h0b ;
            rom[32482] = 8'hfb ;
            rom[32483] = 8'h03 ;
            rom[32484] = 8'h21 ;
            rom[32485] = 8'he6 ;
            rom[32486] = 8'hfc ;
            rom[32487] = 8'hc3 ;
            rom[32488] = 8'h0a ;
            rom[32489] = 8'h11 ;
            rom[32490] = 8'hf4 ;
            rom[32491] = 8'h05 ;
            rom[32492] = 8'hee ;
            rom[32493] = 8'h0a ;
            rom[32494] = 8'hef ;
            rom[32495] = 8'hff ;
            rom[32496] = 8'hd5 ;
            rom[32497] = 8'hea ;
            rom[32498] = 8'h0f ;
            rom[32499] = 8'hf7 ;
            rom[32500] = 8'hff ;
            rom[32501] = 8'h11 ;
            rom[32502] = 8'h1b ;
            rom[32503] = 8'h1c ;
            rom[32504] = 8'h16 ;
            rom[32505] = 8'h07 ;
            rom[32506] = 8'hd7 ;
            rom[32507] = 8'h08 ;
            rom[32508] = 8'hf9 ;
            rom[32509] = 8'h07 ;
            rom[32510] = 8'h1a ;
            rom[32511] = 8'h04 ;
            rom[32512] = 8'he8 ;
            rom[32513] = 8'he9 ;
            rom[32514] = 8'hf4 ;
            rom[32515] = 8'hff ;
            rom[32516] = 8'h05 ;
            rom[32517] = 8'he2 ;
            rom[32518] = 8'h0d ;
            rom[32519] = 8'hfa ;
            rom[32520] = 8'he4 ;
            rom[32521] = 8'h15 ;
            rom[32522] = 8'hfe ;
            rom[32523] = 8'h1b ;
            rom[32524] = 8'h0a ;
            rom[32525] = 8'h02 ;
            rom[32526] = 8'he1 ;
            rom[32527] = 8'h08 ;
            rom[32528] = 8'hfa ;
            rom[32529] = 8'h07 ;
            rom[32530] = 8'hde ;
            rom[32531] = 8'hda ;
            rom[32532] = 8'h06 ;
            rom[32533] = 8'h1e ;
            rom[32534] = 8'h08 ;
            rom[32535] = 8'h1d ;
            rom[32536] = 8'hff ;
            rom[32537] = 8'h1c ;
            rom[32538] = 8'h0a ;
            rom[32539] = 8'h01 ;
            rom[32540] = 8'hd1 ;
            rom[32541] = 8'hf6 ;
            rom[32542] = 8'hf1 ;
            rom[32543] = 8'hd8 ;
            rom[32544] = 8'h07 ;
            rom[32545] = 8'h23 ;
            rom[32546] = 8'hf1 ;
            rom[32547] = 8'h04 ;
            rom[32548] = 8'h0f ;
            rom[32549] = 8'h11 ;
            rom[32550] = 8'h02 ;
            rom[32551] = 8'he6 ;
            rom[32552] = 8'hfe ;
            rom[32553] = 8'hce ;
            rom[32554] = 8'hf1 ;
            rom[32555] = 8'hfb ;
            rom[32556] = 8'h13 ;
            rom[32557] = 8'hfa ;
            rom[32558] = 8'h01 ;
            rom[32559] = 8'hca ;
            rom[32560] = 8'hd6 ;
            rom[32561] = 8'hec ;
            rom[32562] = 8'he6 ;
            rom[32563] = 8'hf4 ;
            rom[32564] = 8'h11 ;
            rom[32565] = 8'hd2 ;
            rom[32566] = 8'hf7 ;
            rom[32567] = 8'hd6 ;
            rom[32568] = 8'hf0 ;
            rom[32569] = 8'h0c ;
            rom[32570] = 8'hfd ;
            rom[32571] = 8'h16 ;
            rom[32572] = 8'hf9 ;
            rom[32573] = 8'hd5 ;
            rom[32574] = 8'h00 ;
            rom[32575] = 8'hff ;
            rom[32576] = 8'hfa ;
            rom[32577] = 8'hff ;
            rom[32578] = 8'he4 ;
            rom[32579] = 8'hdd ;
            rom[32580] = 8'hd4 ;
            rom[32581] = 8'hfa ;
            rom[32582] = 8'hbb ;
            rom[32583] = 8'h08 ;
            rom[32584] = 8'hde ;
            rom[32585] = 8'hef ;
            rom[32586] = 8'h39 ;
            rom[32587] = 8'h1e ;
            rom[32588] = 8'hf9 ;
            rom[32589] = 8'h00 ;
            rom[32590] = 8'hff ;
            rom[32591] = 8'h22 ;
            rom[32592] = 8'hd9 ;
            rom[32593] = 8'hfc ;
            rom[32594] = 8'h07 ;
            rom[32595] = 8'h09 ;
            rom[32596] = 8'h05 ;
            rom[32597] = 8'he7 ;
            rom[32598] = 8'hd6 ;
            rom[32599] = 8'h09 ;
            rom[32600] = 8'h2b ;
            rom[32601] = 8'h0a ;
            rom[32602] = 8'he5 ;
            rom[32603] = 8'h0b ;
            rom[32604] = 8'h16 ;
            rom[32605] = 8'hf7 ;
            rom[32606] = 8'h02 ;
            rom[32607] = 8'h1a ;
            rom[32608] = 8'h10 ;
            rom[32609] = 8'hed ;
            rom[32610] = 8'h10 ;
            rom[32611] = 8'hec ;
            rom[32612] = 8'h13 ;
            rom[32613] = 8'h06 ;
            rom[32614] = 8'hf7 ;
            rom[32615] = 8'h09 ;
            rom[32616] = 8'hf1 ;
            rom[32617] = 8'h06 ;
            rom[32618] = 8'hda ;
            rom[32619] = 8'h11 ;
            rom[32620] = 8'h00 ;
            rom[32621] = 8'h0d ;
            rom[32622] = 8'h0d ;
            rom[32623] = 8'h29 ;
            rom[32624] = 8'h1a ;
            rom[32625] = 8'h05 ;
            rom[32626] = 8'h0c ;
            rom[32627] = 8'h0a ;
            rom[32628] = 8'h02 ;
            rom[32629] = 8'hfc ;
            rom[32630] = 8'h0b ;
            rom[32631] = 8'h0a ;
            rom[32632] = 8'h0e ;
            rom[32633] = 8'hff ;
            rom[32634] = 8'h13 ;
            rom[32635] = 8'hdc ;
            rom[32636] = 8'hee ;
            rom[32637] = 8'hfa ;
            rom[32638] = 8'hc9 ;
            rom[32639] = 8'hf2 ;
            rom[32640] = 8'hf7 ;
            rom[32641] = 8'h0a ;
            rom[32642] = 8'hdd ;
            rom[32643] = 8'hf0 ;
            rom[32644] = 8'h12 ;
            rom[32645] = 8'hf2 ;
            rom[32646] = 8'he4 ;
            rom[32647] = 8'hf4 ;
            rom[32648] = 8'h0d ;
            rom[32649] = 8'hf8 ;
            rom[32650] = 8'hbd ;
            rom[32651] = 8'he4 ;
            rom[32652] = 8'h1b ;
            rom[32653] = 8'hea ;
            rom[32654] = 8'h12 ;
            rom[32655] = 8'hf9 ;
            rom[32656] = 8'h13 ;
            rom[32657] = 8'hf9 ;
            rom[32658] = 8'h00 ;
            rom[32659] = 8'hf5 ;
            rom[32660] = 8'hc0 ;
            rom[32661] = 8'h06 ;
            rom[32662] = 8'hb7 ;
            rom[32663] = 8'hfe ;
            rom[32664] = 8'hdc ;
            rom[32665] = 8'hfe ;
            rom[32666] = 8'hc2 ;
            rom[32667] = 8'hee ;
            rom[32668] = 8'hfd ;
            rom[32669] = 8'h0f ;
            rom[32670] = 8'hae ;
            rom[32671] = 8'he9 ;
            rom[32672] = 8'h09 ;
            rom[32673] = 8'he7 ;
            rom[32674] = 8'h03 ;
            rom[32675] = 8'hfa ;
            rom[32676] = 8'he5 ;
            rom[32677] = 8'hd7 ;
            rom[32678] = 8'h00 ;
            rom[32679] = 8'he3 ;
            rom[32680] = 8'h03 ;
            rom[32681] = 8'h15 ;
            rom[32682] = 8'h13 ;
            rom[32683] = 8'hff ;
            rom[32684] = 8'h08 ;
            rom[32685] = 8'hfa ;
            rom[32686] = 8'h10 ;
            rom[32687] = 8'heb ;
            rom[32688] = 8'hec ;
            rom[32689] = 8'hfc ;
            rom[32690] = 8'he9 ;
            rom[32691] = 8'h19 ;
            rom[32692] = 8'h01 ;
            rom[32693] = 8'h1c ;
            rom[32694] = 8'hfb ;
            rom[32695] = 8'hf0 ;
            rom[32696] = 8'hf6 ;
            rom[32697] = 8'hfe ;
            rom[32698] = 8'hf7 ;
            rom[32699] = 8'he9 ;
            rom[32700] = 8'h00 ;
            rom[32701] = 8'hcc ;
            rom[32702] = 8'hfa ;
            rom[32703] = 8'h15 ;
            rom[32704] = 8'h16 ;
            rom[32705] = 8'hfa ;
            rom[32706] = 8'he6 ;
            rom[32707] = 8'hf4 ;
            rom[32708] = 8'hde ;
            rom[32709] = 8'h07 ;
            rom[32710] = 8'h0e ;
            rom[32711] = 8'hfc ;
            rom[32712] = 8'he8 ;
            rom[32713] = 8'hef ;
            rom[32714] = 8'hff ;
            rom[32715] = 8'h0f ;
            rom[32716] = 8'h0b ;
            rom[32717] = 8'hce ;
            rom[32718] = 8'h0c ;
            rom[32719] = 8'hef ;
            rom[32720] = 8'h09 ;
            rom[32721] = 8'hd4 ;
            rom[32722] = 8'hfc ;
            rom[32723] = 8'he6 ;
            rom[32724] = 8'h0a ;
            rom[32725] = 8'h10 ;
            rom[32726] = 8'hea ;
            rom[32727] = 8'h0d ;
            rom[32728] = 8'h0a ;
            rom[32729] = 8'hd9 ;
            rom[32730] = 8'h24 ;
            rom[32731] = 8'h05 ;
            rom[32732] = 8'hd6 ;
            rom[32733] = 8'hd1 ;
            rom[32734] = 8'he9 ;
            rom[32735] = 8'hfd ;
            rom[32736] = 8'h04 ;
            rom[32737] = 8'hfd ;
            rom[32738] = 8'h01 ;
            rom[32739] = 8'hfa ;
            rom[32740] = 8'h01 ;
            rom[32741] = 8'h06 ;
            rom[32742] = 8'hfc ;
            rom[32743] = 8'h15 ;
            rom[32744] = 8'he7 ;
            rom[32745] = 8'h06 ;
            rom[32746] = 8'h07 ;
            rom[32747] = 8'hd1 ;
            rom[32748] = 8'hfd ;
            rom[32749] = 8'hdf ;
            rom[32750] = 8'hef ;
            rom[32751] = 8'he5 ;
            rom[32752] = 8'hf5 ;
            rom[32753] = 8'hf5 ;
            rom[32754] = 8'h2c ;
            rom[32755] = 8'he0 ;
            rom[32756] = 8'hfd ;
            rom[32757] = 8'hf9 ;
            rom[32758] = 8'hf2 ;
            rom[32759] = 8'h0c ;
            rom[32760] = 8'h0e ;
            rom[32761] = 8'hbc ;
            rom[32762] = 8'hf0 ;
            rom[32763] = 8'hd0 ;
            rom[32764] = 8'hfd ;
            rom[32765] = 8'he7 ;
            rom[32766] = 8'hf1 ;
            rom[32767] = 8'hf6 ;
            rom[32768] = 8'h19 ;
            rom[32769] = 8'hf6 ;
            rom[32770] = 8'h13 ;
            rom[32771] = 8'hed ;
            rom[32772] = 8'he5 ;
            rom[32773] = 8'h11 ;
            rom[32774] = 8'hfb ;
            rom[32775] = 8'h0f ;
            rom[32776] = 8'heb ;
            rom[32777] = 8'hff ;
            rom[32778] = 8'h06 ;
            rom[32779] = 8'h00 ;
            rom[32780] = 8'h0e ;
            rom[32781] = 8'hf5 ;
            rom[32782] = 8'h37 ;
            rom[32783] = 8'h04 ;
            rom[32784] = 8'hfd ;
            rom[32785] = 8'he9 ;
            rom[32786] = 8'h03 ;
            rom[32787] = 8'hee ;
            rom[32788] = 8'h00 ;
            rom[32789] = 8'h1a ;
            rom[32790] = 8'hfa ;
            rom[32791] = 8'hcf ;
            rom[32792] = 8'hf2 ;
            rom[32793] = 8'hf4 ;
            rom[32794] = 8'hef ;
            rom[32795] = 8'hfc ;
            rom[32796] = 8'h17 ;
            rom[32797] = 8'hf6 ;
            rom[32798] = 8'he5 ;
            rom[32799] = 8'he9 ;
            rom[32800] = 8'hfe ;
            rom[32801] = 8'hef ;
            rom[32802] = 8'hee ;
            rom[32803] = 8'h1a ;
            rom[32804] = 8'h2a ;
            rom[32805] = 8'h05 ;
            rom[32806] = 8'h27 ;
            rom[32807] = 8'hee ;
            rom[32808] = 8'h0c ;
            rom[32809] = 8'hb9 ;
            rom[32810] = 8'h11 ;
            rom[32811] = 8'hdf ;
            rom[32812] = 8'hf5 ;
            rom[32813] = 8'h17 ;
            rom[32814] = 8'h28 ;
            rom[32815] = 8'hf2 ;
            rom[32816] = 8'hd1 ;
            rom[32817] = 8'hff ;
            rom[32818] = 8'h00 ;
            rom[32819] = 8'hd3 ;
            rom[32820] = 8'hec ;
            rom[32821] = 8'h21 ;
            rom[32822] = 8'h05 ;
            rom[32823] = 8'he8 ;
            rom[32824] = 8'h20 ;
            rom[32825] = 8'h11 ;
            rom[32826] = 8'hfc ;
            rom[32827] = 8'hfc ;
            rom[32828] = 8'h09 ;
            rom[32829] = 8'hf1 ;
            rom[32830] = 8'he0 ;
            rom[32831] = 8'he9 ;
            rom[32832] = 8'h06 ;
            rom[32833] = 8'h0c ;
            rom[32834] = 8'hf6 ;
            rom[32835] = 8'hfb ;
            rom[32836] = 8'he4 ;
            rom[32837] = 8'h0b ;
            rom[32838] = 8'h03 ;
            rom[32839] = 8'h23 ;
            rom[32840] = 8'hf2 ;
            rom[32841] = 8'h0f ;
            rom[32842] = 8'hee ;
            rom[32843] = 8'hf9 ;
            rom[32844] = 8'hde ;
            rom[32845] = 8'hf8 ;
            rom[32846] = 8'hed ;
            rom[32847] = 8'he9 ;
            rom[32848] = 8'h03 ;
            rom[32849] = 8'hde ;
            rom[32850] = 8'h05 ;
            rom[32851] = 8'h06 ;
            rom[32852] = 8'h05 ;
            rom[32853] = 8'hcf ;
            rom[32854] = 8'h13 ;
            rom[32855] = 8'hdd ;
            rom[32856] = 8'h09 ;
            rom[32857] = 8'hde ;
            rom[32858] = 8'h14 ;
            rom[32859] = 8'he4 ;
            rom[32860] = 8'he6 ;
            rom[32861] = 8'he1 ;
            rom[32862] = 8'he2 ;
            rom[32863] = 8'hd8 ;
            rom[32864] = 8'hf6 ;
            rom[32865] = 8'h12 ;
            rom[32866] = 8'hff ;
            rom[32867] = 8'hec ;
            rom[32868] = 8'hef ;
            rom[32869] = 8'he3 ;
            rom[32870] = 8'hed ;
            rom[32871] = 8'h03 ;
            rom[32872] = 8'h1a ;
            rom[32873] = 8'h2a ;
            rom[32874] = 8'hdb ;
            rom[32875] = 8'hdf ;
            rom[32876] = 8'h0a ;
            rom[32877] = 8'h2f ;
            rom[32878] = 8'h05 ;
            rom[32879] = 8'hff ;
            rom[32880] = 8'h08 ;
            rom[32881] = 8'hfe ;
            rom[32882] = 8'h18 ;
            rom[32883] = 8'h1d ;
            rom[32884] = 8'h0d ;
            rom[32885] = 8'h11 ;
            rom[32886] = 8'hf5 ;
            rom[32887] = 8'hf6 ;
            rom[32888] = 8'h07 ;
            rom[32889] = 8'h23 ;
            rom[32890] = 8'hfd ;
            rom[32891] = 8'he1 ;
            rom[32892] = 8'h0d ;
            rom[32893] = 8'hda ;
            rom[32894] = 8'hfb ;
            rom[32895] = 8'h0d ;
            rom[32896] = 8'h05 ;
            rom[32897] = 8'h0a ;
            rom[32898] = 8'hda ;
            rom[32899] = 8'h0b ;
            rom[32900] = 8'hfe ;
            rom[32901] = 8'h00 ;
            rom[32902] = 8'hd8 ;
            rom[32903] = 8'h10 ;
            rom[32904] = 8'hfd ;
            rom[32905] = 8'heb ;
            rom[32906] = 8'h03 ;
            rom[32907] = 8'he4 ;
            rom[32908] = 8'hda ;
            rom[32909] = 8'h01 ;
            rom[32910] = 8'h1a ;
            rom[32911] = 8'hfd ;
            rom[32912] = 8'he0 ;
            rom[32913] = 8'h01 ;
            rom[32914] = 8'he5 ;
            rom[32915] = 8'h12 ;
            rom[32916] = 8'he7 ;
            rom[32917] = 8'hf4 ;
            rom[32918] = 8'hea ;
            rom[32919] = 8'hfa ;
            rom[32920] = 8'h02 ;
            rom[32921] = 8'hfc ;
            rom[32922] = 8'h10 ;
            rom[32923] = 8'hf1 ;
            rom[32924] = 8'h06 ;
            rom[32925] = 8'hdb ;
            rom[32926] = 8'h06 ;
            rom[32927] = 8'hf0 ;
            rom[32928] = 8'he3 ;
            rom[32929] = 8'h12 ;
            rom[32930] = 8'hf7 ;
            rom[32931] = 8'hf9 ;
            rom[32932] = 8'hcf ;
            rom[32933] = 8'he5 ;
            rom[32934] = 8'hea ;
            rom[32935] = 8'hfc ;
            rom[32936] = 8'h02 ;
            rom[32937] = 8'he0 ;
            rom[32938] = 8'h13 ;
            rom[32939] = 8'hdc ;
            rom[32940] = 8'h05 ;
            rom[32941] = 8'he1 ;
            rom[32942] = 8'h05 ;
            rom[32943] = 8'hff ;
            rom[32944] = 8'hd7 ;
            rom[32945] = 8'hfe ;
            rom[32946] = 8'hfa ;
            rom[32947] = 8'h0c ;
            rom[32948] = 8'h17 ;
            rom[32949] = 8'he3 ;
            rom[32950] = 8'hdd ;
            rom[32951] = 8'hfc ;
            rom[32952] = 8'h0c ;
            rom[32953] = 8'hf9 ;
            rom[32954] = 8'hfb ;
            rom[32955] = 8'he5 ;
            rom[32956] = 8'hdf ;
            rom[32957] = 8'h0b ;
            rom[32958] = 8'hbd ;
            rom[32959] = 8'hfb ;
            rom[32960] = 8'h02 ;
            rom[32961] = 8'he0 ;
            rom[32962] = 8'h07 ;
            rom[32963] = 8'hd9 ;
            rom[32964] = 8'h0a ;
            rom[32965] = 8'hd1 ;
            rom[32966] = 8'hff ;
            rom[32967] = 8'hb9 ;
            rom[32968] = 8'h02 ;
            rom[32969] = 8'hd2 ;
            rom[32970] = 8'h10 ;
            rom[32971] = 8'hfa ;
            rom[32972] = 8'he8 ;
            rom[32973] = 8'h16 ;
            rom[32974] = 8'h05 ;
            rom[32975] = 8'hfe ;
            rom[32976] = 8'heb ;
            rom[32977] = 8'h02 ;
            rom[32978] = 8'hc3 ;
            rom[32979] = 8'hf8 ;
            rom[32980] = 8'h0d ;
            rom[32981] = 8'he1 ;
            rom[32982] = 8'hf0 ;
            rom[32983] = 8'hdc ;
            rom[32984] = 8'hfe ;
            rom[32985] = 8'hfe ;
            rom[32986] = 8'hd6 ;
            rom[32987] = 8'hec ;
            rom[32988] = 8'hed ;
            rom[32989] = 8'hfd ;
            rom[32990] = 8'hf6 ;
            rom[32991] = 8'he9 ;
            rom[32992] = 8'hf2 ;
            rom[32993] = 8'hf0 ;
            rom[32994] = 8'hdd ;
            rom[32995] = 8'hcd ;
            rom[32996] = 8'heb ;
            rom[32997] = 8'hd2 ;
            rom[32998] = 8'hd3 ;
            rom[32999] = 8'hea ;
            rom[33000] = 8'heb ;
            rom[33001] = 8'hc3 ;
            rom[33002] = 8'hdc ;
            rom[33003] = 8'h02 ;
            rom[33004] = 8'hf7 ;
            rom[33005] = 8'hd9 ;
            rom[33006] = 8'hf8 ;
            rom[33007] = 8'h00 ;
            rom[33008] = 8'hed ;
            rom[33009] = 8'hfc ;
            rom[33010] = 8'h16 ;
            rom[33011] = 8'hed ;
            rom[33012] = 8'h07 ;
            rom[33013] = 8'hf3 ;
            rom[33014] = 8'h03 ;
            rom[33015] = 8'he1 ;
            rom[33016] = 8'hdb ;
            rom[33017] = 8'h12 ;
            rom[33018] = 8'h08 ;
            rom[33019] = 8'hf8 ;
            rom[33020] = 8'h08 ;
            rom[33021] = 8'hca ;
            rom[33022] = 8'hdc ;
            rom[33023] = 8'he5 ;
            rom[33024] = 8'h11 ;
            rom[33025] = 8'hf6 ;
            rom[33026] = 8'hde ;
            rom[33027] = 8'h0f ;
            rom[33028] = 8'hf8 ;
            rom[33029] = 8'hd1 ;
            rom[33030] = 8'h08 ;
            rom[33031] = 8'hdc ;
            rom[33032] = 8'h0a ;
            rom[33033] = 8'h1f ;
            rom[33034] = 8'hec ;
            rom[33035] = 8'he2 ;
            rom[33036] = 8'he0 ;
            rom[33037] = 8'hb3 ;
            rom[33038] = 8'h04 ;
            rom[33039] = 8'hfe ;
            rom[33040] = 8'hf7 ;
            rom[33041] = 8'hf2 ;
            rom[33042] = 8'h27 ;
            rom[33043] = 8'h00 ;
            rom[33044] = 8'hec ;
            rom[33045] = 8'h17 ;
            rom[33046] = 8'hdc ;
            rom[33047] = 8'hf0 ;
            rom[33048] = 8'h0c ;
            rom[33049] = 8'hf7 ;
            rom[33050] = 8'h01 ;
            rom[33051] = 8'h0b ;
            rom[33052] = 8'hc5 ;
            rom[33053] = 8'h28 ;
            rom[33054] = 8'hfa ;
            rom[33055] = 8'hf3 ;
            rom[33056] = 8'hef ;
            rom[33057] = 8'heb ;
            rom[33058] = 8'h11 ;
            rom[33059] = 8'hff ;
            rom[33060] = 8'h02 ;
            rom[33061] = 8'h06 ;
            rom[33062] = 8'hc3 ;
            rom[33063] = 8'hcc ;
            rom[33064] = 8'hee ;
            rom[33065] = 8'h00 ;
            rom[33066] = 8'h0e ;
            rom[33067] = 8'hf2 ;
            rom[33068] = 8'h1c ;
            rom[33069] = 8'h0d ;
            rom[33070] = 8'h19 ;
            rom[33071] = 8'h0a ;
            rom[33072] = 8'h0f ;
            rom[33073] = 8'h04 ;
            rom[33074] = 8'hde ;
            rom[33075] = 8'hde ;
            rom[33076] = 8'h1b ;
            rom[33077] = 8'hd3 ;
            rom[33078] = 8'hdc ;
            rom[33079] = 8'hf6 ;
            rom[33080] = 8'h1c ;
            rom[33081] = 8'h1f ;
            rom[33082] = 8'h12 ;
            rom[33083] = 8'hea ;
            rom[33084] = 8'hf5 ;
            rom[33085] = 8'hc8 ;
            rom[33086] = 8'he3 ;
            rom[33087] = 8'h00 ;
            rom[33088] = 8'hf2 ;
            rom[33089] = 8'h15 ;
            rom[33090] = 8'h15 ;
            rom[33091] = 8'h0d ;
            rom[33092] = 8'hf7 ;
            rom[33093] = 8'h06 ;
            rom[33094] = 8'hd2 ;
            rom[33095] = 8'h12 ;
            rom[33096] = 8'hed ;
            rom[33097] = 8'hfe ;
            rom[33098] = 8'h13 ;
            rom[33099] = 8'he6 ;
            rom[33100] = 8'hfe ;
            rom[33101] = 8'hff ;
            rom[33102] = 8'he5 ;
            rom[33103] = 8'h0c ;
            rom[33104] = 8'h0d ;
            rom[33105] = 8'hc1 ;
            rom[33106] = 8'hfd ;
            rom[33107] = 8'hf4 ;
            rom[33108] = 8'he4 ;
            rom[33109] = 8'h06 ;
            rom[33110] = 8'hc6 ;
            rom[33111] = 8'h0e ;
            rom[33112] = 8'h24 ;
            rom[33113] = 8'hf0 ;
            rom[33114] = 8'h10 ;
            rom[33115] = 8'hfc ;
            rom[33116] = 8'he5 ;
            rom[33117] = 8'hd8 ;
            rom[33118] = 8'hfc ;
            rom[33119] = 8'h1f ;
            rom[33120] = 8'hf4 ;
            rom[33121] = 8'hd2 ;
            rom[33122] = 8'hff ;
            rom[33123] = 8'h0e ;
            rom[33124] = 8'heb ;
            rom[33125] = 8'h12 ;
            rom[33126] = 8'h0c ;
            rom[33127] = 8'h07 ;
            rom[33128] = 8'hdf ;
            rom[33129] = 8'hcc ;
            rom[33130] = 8'h06 ;
            rom[33131] = 8'h16 ;
            rom[33132] = 8'hfa ;
            rom[33133] = 8'hf6 ;
            rom[33134] = 8'hfc ;
            rom[33135] = 8'h05 ;
            rom[33136] = 8'h11 ;
            rom[33137] = 8'h14 ;
            rom[33138] = 8'h03 ;
            rom[33139] = 8'hf2 ;
            rom[33140] = 8'hec ;
            rom[33141] = 8'h07 ;
            rom[33142] = 8'h02 ;
            rom[33143] = 8'h16 ;
            rom[33144] = 8'hf2 ;
            rom[33145] = 8'h13 ;
            rom[33146] = 8'he6 ;
            rom[33147] = 8'hf9 ;
            rom[33148] = 8'hff ;
            rom[33149] = 8'hf8 ;
            rom[33150] = 8'heb ;
            rom[33151] = 8'heb ;
            rom[33152] = 8'hba ;
            rom[33153] = 8'h02 ;
            rom[33154] = 8'h14 ;
            rom[33155] = 8'hfc ;
            rom[33156] = 8'hec ;
            rom[33157] = 8'h08 ;
            rom[33158] = 8'h1d ;
            rom[33159] = 8'h00 ;
            rom[33160] = 8'hf2 ;
            rom[33161] = 8'h0a ;
            rom[33162] = 8'hc5 ;
            rom[33163] = 8'h03 ;
            rom[33164] = 8'h10 ;
            rom[33165] = 8'he3 ;
            rom[33166] = 8'h04 ;
            rom[33167] = 8'hf8 ;
            rom[33168] = 8'h00 ;
            rom[33169] = 8'hc8 ;
            rom[33170] = 8'hff ;
            rom[33171] = 8'hd4 ;
            rom[33172] = 8'h07 ;
            rom[33173] = 8'hf5 ;
            rom[33174] = 8'h00 ;
            rom[33175] = 8'he1 ;
            rom[33176] = 8'hf3 ;
            rom[33177] = 8'h09 ;
            rom[33178] = 8'hff ;
            rom[33179] = 8'hf0 ;
            rom[33180] = 8'h04 ;
            rom[33181] = 8'h13 ;
            rom[33182] = 8'h03 ;
            rom[33183] = 8'hea ;
            rom[33184] = 8'h00 ;
            rom[33185] = 8'hd5 ;
            rom[33186] = 8'hd5 ;
            rom[33187] = 8'h0a ;
            rom[33188] = 8'h04 ;
            rom[33189] = 8'hf7 ;
            rom[33190] = 8'h0c ;
            rom[33191] = 8'h02 ;
            rom[33192] = 8'h0b ;
            rom[33193] = 8'hdb ;
            rom[33194] = 8'h18 ;
            rom[33195] = 8'hf9 ;
            rom[33196] = 8'h14 ;
            rom[33197] = 8'he5 ;
            rom[33198] = 8'hfb ;
            rom[33199] = 8'hfa ;
            rom[33200] = 8'h0a ;
            rom[33201] = 8'h04 ;
            rom[33202] = 8'h05 ;
            rom[33203] = 8'hfb ;
            rom[33204] = 8'hec ;
            rom[33205] = 8'h22 ;
            rom[33206] = 8'h00 ;
            rom[33207] = 8'he7 ;
            rom[33208] = 8'hfb ;
            rom[33209] = 8'hfe ;
            rom[33210] = 8'h02 ;
            rom[33211] = 8'hf6 ;
            rom[33212] = 8'h09 ;
            rom[33213] = 8'hff ;
            rom[33214] = 8'hf4 ;
            rom[33215] = 8'he4 ;
            rom[33216] = 8'h07 ;
            rom[33217] = 8'hed ;
            rom[33218] = 8'hfc ;
            rom[33219] = 8'hfc ;
            rom[33220] = 8'he2 ;
            rom[33221] = 8'h03 ;
            rom[33222] = 8'hfa ;
            rom[33223] = 8'h0f ;
            rom[33224] = 8'hb3 ;
            rom[33225] = 8'hf7 ;
            rom[33226] = 8'h17 ;
            rom[33227] = 8'h13 ;
            rom[33228] = 8'hff ;
            rom[33229] = 8'he8 ;
            rom[33230] = 8'hd3 ;
            rom[33231] = 8'he6 ;
            rom[33232] = 8'h02 ;
            rom[33233] = 8'he7 ;
            rom[33234] = 8'h04 ;
            rom[33235] = 8'h00 ;
            rom[33236] = 8'hd2 ;
            rom[33237] = 8'h0d ;
            rom[33238] = 8'hee ;
            rom[33239] = 8'hdb ;
            rom[33240] = 8'hf9 ;
            rom[33241] = 8'h18 ;
            rom[33242] = 8'h18 ;
            rom[33243] = 8'h00 ;
            rom[33244] = 8'hed ;
            rom[33245] = 8'hdb ;
            rom[33246] = 8'hec ;
            rom[33247] = 8'hfb ;
            rom[33248] = 8'h07 ;
            rom[33249] = 8'h0b ;
            rom[33250] = 8'hf9 ;
            rom[33251] = 8'hf7 ;
            rom[33252] = 8'h28 ;
            rom[33253] = 8'hf1 ;
            rom[33254] = 8'hfc ;
            rom[33255] = 8'he9 ;
            rom[33256] = 8'h14 ;
            rom[33257] = 8'hdd ;
            rom[33258] = 8'hfb ;
            rom[33259] = 8'h0e ;
            rom[33260] = 8'hfa ;
            rom[33261] = 8'h16 ;
            rom[33262] = 8'hb3 ;
            rom[33263] = 8'h13 ;
            rom[33264] = 8'h09 ;
            rom[33265] = 8'hf9 ;
            rom[33266] = 8'h05 ;
            rom[33267] = 8'hff ;
            rom[33268] = 8'he2 ;
            rom[33269] = 8'h17 ;
            rom[33270] = 8'hff ;
            rom[33271] = 8'hfb ;
            rom[33272] = 8'hf5 ;
            rom[33273] = 8'hdc ;
            rom[33274] = 8'h0c ;
            rom[33275] = 8'h24 ;
            rom[33276] = 8'hed ;
            rom[33277] = 8'he0 ;
            rom[33278] = 8'hf3 ;
            rom[33279] = 8'h11 ;
            rom[33280] = 8'h0a ;
            rom[33281] = 8'h0e ;
            rom[33282] = 8'h30 ;
            rom[33283] = 8'h0c ;
            rom[33284] = 8'h1e ;
            rom[33285] = 8'hc6 ;
            rom[33286] = 8'hfb ;
            rom[33287] = 8'hf9 ;
            rom[33288] = 8'h1a ;
            rom[33289] = 8'h01 ;
            rom[33290] = 8'hd8 ;
            rom[33291] = 8'hf1 ;
            rom[33292] = 8'he3 ;
            rom[33293] = 8'h0a ;
            rom[33294] = 8'hdd ;
            rom[33295] = 8'he3 ;
            rom[33296] = 8'h13 ;
            rom[33297] = 8'hfe ;
            rom[33298] = 8'h32 ;
            rom[33299] = 8'heb ;
            rom[33300] = 8'h0e ;
            rom[33301] = 8'h21 ;
            rom[33302] = 8'h10 ;
            rom[33303] = 8'hf9 ;
            rom[33304] = 8'h06 ;
            rom[33305] = 8'h0f ;
            rom[33306] = 8'he4 ;
            rom[33307] = 8'h1f ;
            rom[33308] = 8'h07 ;
            rom[33309] = 8'hf1 ;
            rom[33310] = 8'h33 ;
            rom[33311] = 8'h07 ;
            rom[33312] = 8'hf0 ;
            rom[33313] = 8'h21 ;
            rom[33314] = 8'h0a ;
            rom[33315] = 8'hc0 ;
            rom[33316] = 8'h1d ;
            rom[33317] = 8'h04 ;
            rom[33318] = 8'hff ;
            rom[33319] = 8'h06 ;
            rom[33320] = 8'hea ;
            rom[33321] = 8'h06 ;
            rom[33322] = 8'he1 ;
            rom[33323] = 8'hdf ;
            rom[33324] = 8'hfc ;
            rom[33325] = 8'hfb ;
            rom[33326] = 8'hdd ;
            rom[33327] = 8'h23 ;
            rom[33328] = 8'hec ;
            rom[33329] = 8'h16 ;
            rom[33330] = 8'hed ;
            rom[33331] = 8'hfb ;
            rom[33332] = 8'he4 ;
            rom[33333] = 8'he6 ;
            rom[33334] = 8'he6 ;
            rom[33335] = 8'hfe ;
            rom[33336] = 8'he8 ;
            rom[33337] = 8'hf5 ;
            rom[33338] = 8'hf1 ;
            rom[33339] = 8'h09 ;
            rom[33340] = 8'h1b ;
            rom[33341] = 8'h09 ;
            rom[33342] = 8'hc4 ;
            rom[33343] = 8'hf3 ;
            rom[33344] = 8'hea ;
            rom[33345] = 8'hfd ;
            rom[33346] = 8'hfa ;
            rom[33347] = 8'hff ;
            rom[33348] = 8'h29 ;
            rom[33349] = 8'h01 ;
            rom[33350] = 8'hf2 ;
            rom[33351] = 8'h00 ;
            rom[33352] = 8'h0f ;
            rom[33353] = 8'hf6 ;
            rom[33354] = 8'hfd ;
            rom[33355] = 8'h07 ;
            rom[33356] = 8'h01 ;
            rom[33357] = 8'hdd ;
            rom[33358] = 8'haf ;
            rom[33359] = 8'hf8 ;
            rom[33360] = 8'hf2 ;
            rom[33361] = 8'h1f ;
            rom[33362] = 8'hd0 ;
            rom[33363] = 8'h0b ;
            rom[33364] = 8'h0c ;
            rom[33365] = 8'hd3 ;
            rom[33366] = 8'h13 ;
            rom[33367] = 8'h0c ;
            rom[33368] = 8'hf7 ;
            rom[33369] = 8'h11 ;
            rom[33370] = 8'hfb ;
            rom[33371] = 8'ha6 ;
            rom[33372] = 8'h00 ;
            rom[33373] = 8'h00 ;
            rom[33374] = 8'hf4 ;
            rom[33375] = 8'hc7 ;
            rom[33376] = 8'h0f ;
            rom[33377] = 8'h0f ;
            rom[33378] = 8'he8 ;
            rom[33379] = 8'hed ;
            rom[33380] = 8'he7 ;
            rom[33381] = 8'he0 ;
            rom[33382] = 8'h13 ;
            rom[33383] = 8'hef ;
            rom[33384] = 8'hf9 ;
            rom[33385] = 8'h13 ;
            rom[33386] = 8'h11 ;
            rom[33387] = 8'hd5 ;
            rom[33388] = 8'hba ;
            rom[33389] = 8'hec ;
            rom[33390] = 8'hf1 ;
            rom[33391] = 8'h11 ;
            rom[33392] = 8'he3 ;
            rom[33393] = 8'h06 ;
            rom[33394] = 8'hf4 ;
            rom[33395] = 8'hf4 ;
            rom[33396] = 8'hf0 ;
            rom[33397] = 8'hfa ;
            rom[33398] = 8'hfa ;
            rom[33399] = 8'he3 ;
            rom[33400] = 8'hff ;
            rom[33401] = 8'h02 ;
            rom[33402] = 8'hc8 ;
            rom[33403] = 8'h1c ;
            rom[33404] = 8'hd6 ;
            rom[33405] = 8'h18 ;
            rom[33406] = 8'h07 ;
            rom[33407] = 8'hef ;
            rom[33408] = 8'hf5 ;
            rom[33409] = 8'hde ;
            rom[33410] = 8'he3 ;
            rom[33411] = 8'h0a ;
            rom[33412] = 8'h19 ;
            rom[33413] = 8'hf7 ;
            rom[33414] = 8'hf3 ;
            rom[33415] = 8'hfe ;
            rom[33416] = 8'hfd ;
            rom[33417] = 8'h02 ;
            rom[33418] = 8'h1c ;
            rom[33419] = 8'hd6 ;
            rom[33420] = 8'hf4 ;
            rom[33421] = 8'he2 ;
            rom[33422] = 8'h1b ;
            rom[33423] = 8'hf5 ;
            rom[33424] = 8'hed ;
            rom[33425] = 8'heb ;
            rom[33426] = 8'h09 ;
            rom[33427] = 8'hfa ;
            rom[33428] = 8'h0b ;
            rom[33429] = 8'h18 ;
            rom[33430] = 8'hfb ;
            rom[33431] = 8'h07 ;
            rom[33432] = 8'h10 ;
            rom[33433] = 8'h15 ;
            rom[33434] = 8'h1e ;
            rom[33435] = 8'h0d ;
            rom[33436] = 8'hee ;
            rom[33437] = 8'h19 ;
            rom[33438] = 8'h1d ;
            rom[33439] = 8'h13 ;
            rom[33440] = 8'h17 ;
            rom[33441] = 8'hd1 ;
            rom[33442] = 8'hc7 ;
            rom[33443] = 8'hff ;
            rom[33444] = 8'hfb ;
            rom[33445] = 8'hec ;
            rom[33446] = 8'hf3 ;
            rom[33447] = 8'h00 ;
            rom[33448] = 8'h01 ;
            rom[33449] = 8'hf8 ;
            rom[33450] = 8'hfd ;
            rom[33451] = 8'hf5 ;
            rom[33452] = 8'h09 ;
            rom[33453] = 8'h19 ;
            rom[33454] = 8'h07 ;
            rom[33455] = 8'he1 ;
            rom[33456] = 8'hba ;
            rom[33457] = 8'h10 ;
            rom[33458] = 8'h26 ;
            rom[33459] = 8'hed ;
            rom[33460] = 8'h0a ;
            rom[33461] = 8'hfc ;
            rom[33462] = 8'h14 ;
            rom[33463] = 8'hd8 ;
            rom[33464] = 8'hea ;
            rom[33465] = 8'h09 ;
            rom[33466] = 8'h13 ;
            rom[33467] = 8'hd8 ;
            rom[33468] = 8'hfe ;
            rom[33469] = 8'hd9 ;
            rom[33470] = 8'hfd ;
            rom[33471] = 8'hfd ;
            rom[33472] = 8'h0a ;
            rom[33473] = 8'hdb ;
            rom[33474] = 8'h0b ;
            rom[33475] = 8'hf0 ;
            rom[33476] = 8'h11 ;
            rom[33477] = 8'h0a ;
            rom[33478] = 8'hcf ;
            rom[33479] = 8'hf9 ;
            rom[33480] = 8'hee ;
            rom[33481] = 8'h07 ;
            rom[33482] = 8'hf7 ;
            rom[33483] = 8'h0f ;
            rom[33484] = 8'hfe ;
            rom[33485] = 8'hf2 ;
            rom[33486] = 8'hff ;
            rom[33487] = 8'h02 ;
            rom[33488] = 8'hfe ;
            rom[33489] = 8'he8 ;
            rom[33490] = 8'h0c ;
            rom[33491] = 8'he7 ;
            rom[33492] = 8'hed ;
            rom[33493] = 8'h20 ;
            rom[33494] = 8'hfd ;
            rom[33495] = 8'hdf ;
            rom[33496] = 8'hea ;
            rom[33497] = 8'h1d ;
            rom[33498] = 8'hfb ;
            rom[33499] = 8'h06 ;
            rom[33500] = 8'h1a ;
            rom[33501] = 8'h0b ;
            rom[33502] = 8'h0d ;
            rom[33503] = 8'hdf ;
            rom[33504] = 8'he8 ;
            rom[33505] = 8'h0e ;
            rom[33506] = 8'h13 ;
            rom[33507] = 8'hd1 ;
            rom[33508] = 8'h01 ;
            rom[33509] = 8'hff ;
            rom[33510] = 8'hea ;
            rom[33511] = 8'he3 ;
            rom[33512] = 8'h07 ;
            rom[33513] = 8'h02 ;
            rom[33514] = 8'hf4 ;
            rom[33515] = 8'h23 ;
            rom[33516] = 8'h08 ;
            rom[33517] = 8'h0c ;
            rom[33518] = 8'he9 ;
            rom[33519] = 8'h1b ;
            rom[33520] = 8'hf6 ;
            rom[33521] = 8'hfa ;
            rom[33522] = 8'h17 ;
            rom[33523] = 8'hfb ;
            rom[33524] = 8'h0e ;
            rom[33525] = 8'hf2 ;
            rom[33526] = 8'h05 ;
            rom[33527] = 8'hfd ;
            rom[33528] = 8'hb2 ;
            rom[33529] = 8'hf6 ;
            rom[33530] = 8'h15 ;
            rom[33531] = 8'hfd ;
            rom[33532] = 8'hf7 ;
            rom[33533] = 8'hf2 ;
            rom[33534] = 8'hd7 ;
            rom[33535] = 8'hf6 ;
            rom[33536] = 8'hff ;
            rom[33537] = 8'h1d ;
            rom[33538] = 8'h06 ;
            rom[33539] = 8'h13 ;
            rom[33540] = 8'hcc ;
            rom[33541] = 8'hf8 ;
            rom[33542] = 8'hfa ;
            rom[33543] = 8'h0b ;
            rom[33544] = 8'h1d ;
            rom[33545] = 8'ha6 ;
            rom[33546] = 8'hef ;
            rom[33547] = 8'h04 ;
            rom[33548] = 8'hea ;
            rom[33549] = 8'h0f ;
            rom[33550] = 8'h0d ;
            rom[33551] = 8'hf1 ;
            rom[33552] = 8'h07 ;
            rom[33553] = 8'hf0 ;
            rom[33554] = 8'h05 ;
            rom[33555] = 8'hf2 ;
            rom[33556] = 8'hfb ;
            rom[33557] = 8'hfc ;
            rom[33558] = 8'he3 ;
            rom[33559] = 8'h05 ;
            rom[33560] = 8'h0f ;
            rom[33561] = 8'hbf ;
            rom[33562] = 8'h06 ;
            rom[33563] = 8'hcf ;
            rom[33564] = 8'he0 ;
            rom[33565] = 8'h20 ;
            rom[33566] = 8'hc0 ;
            rom[33567] = 8'h05 ;
            rom[33568] = 8'h00 ;
            rom[33569] = 8'he4 ;
            rom[33570] = 8'h07 ;
            rom[33571] = 8'he8 ;
            rom[33572] = 8'h02 ;
            rom[33573] = 8'h14 ;
            rom[33574] = 8'h09 ;
            rom[33575] = 8'hcb ;
            rom[33576] = 8'he1 ;
            rom[33577] = 8'hff ;
            rom[33578] = 8'hee ;
            rom[33579] = 8'h04 ;
            rom[33580] = 8'he9 ;
            rom[33581] = 8'h14 ;
            rom[33582] = 8'hdf ;
            rom[33583] = 8'h02 ;
            rom[33584] = 8'h09 ;
            rom[33585] = 8'h16 ;
            rom[33586] = 8'h02 ;
            rom[33587] = 8'hf2 ;
            rom[33588] = 8'he8 ;
            rom[33589] = 8'hed ;
            rom[33590] = 8'hea ;
            rom[33591] = 8'h07 ;
            rom[33592] = 8'h03 ;
            rom[33593] = 8'hcf ;
            rom[33594] = 8'heb ;
            rom[33595] = 8'he3 ;
            rom[33596] = 8'h11 ;
            rom[33597] = 8'hf9 ;
            rom[33598] = 8'h05 ;
            rom[33599] = 8'hd5 ;
            rom[33600] = 8'h18 ;
            rom[33601] = 8'h0b ;
            rom[33602] = 8'hdd ;
            rom[33603] = 8'hf1 ;
            rom[33604] = 8'h07 ;
            rom[33605] = 8'h18 ;
            rom[33606] = 8'hdf ;
            rom[33607] = 8'hfb ;
            rom[33608] = 8'hf0 ;
            rom[33609] = 8'he5 ;
            rom[33610] = 8'hb9 ;
            rom[33611] = 8'h06 ;
            rom[33612] = 8'hbe ;
            rom[33613] = 8'hf2 ;
            rom[33614] = 8'hfc ;
            rom[33615] = 8'h11 ;
            rom[33616] = 8'hf6 ;
            rom[33617] = 8'h0e ;
            rom[33618] = 8'hdd ;
            rom[33619] = 8'hfe ;
            rom[33620] = 8'hf8 ;
            rom[33621] = 8'hd5 ;
            rom[33622] = 8'hef ;
            rom[33623] = 8'h0b ;
            rom[33624] = 8'hfc ;
            rom[33625] = 8'hed ;
            rom[33626] = 8'hf7 ;
            rom[33627] = 8'h01 ;
            rom[33628] = 8'he8 ;
            rom[33629] = 8'h05 ;
            rom[33630] = 8'hf8 ;
            rom[33631] = 8'h09 ;
            rom[33632] = 8'hfd ;
            rom[33633] = 8'h04 ;
            rom[33634] = 8'hf4 ;
            rom[33635] = 8'h1b ;
            rom[33636] = 8'hcb ;
            rom[33637] = 8'h09 ;
            rom[33638] = 8'hef ;
            rom[33639] = 8'hdf ;
            rom[33640] = 8'h1e ;
            rom[33641] = 8'h0c ;
            rom[33642] = 8'h01 ;
            rom[33643] = 8'hfd ;
            rom[33644] = 8'hf8 ;
            rom[33645] = 8'h05 ;
            rom[33646] = 8'h12 ;
            rom[33647] = 8'hd8 ;
            rom[33648] = 8'hf9 ;
            rom[33649] = 8'h18 ;
            rom[33650] = 8'h01 ;
            rom[33651] = 8'h04 ;
            rom[33652] = 8'he9 ;
            rom[33653] = 8'hf8 ;
            rom[33654] = 8'hf8 ;
            rom[33655] = 8'hfb ;
            rom[33656] = 8'he1 ;
            rom[33657] = 8'hee ;
            rom[33658] = 8'ha5 ;
            rom[33659] = 8'h00 ;
            rom[33660] = 8'hf4 ;
            rom[33661] = 8'h10 ;
            rom[33662] = 8'hf9 ;
            rom[33663] = 8'hec ;
            rom[33664] = 8'hf7 ;
            rom[33665] = 8'hd9 ;
            rom[33666] = 8'he8 ;
            rom[33667] = 8'h0b ;
            rom[33668] = 8'hd2 ;
            rom[33669] = 8'he4 ;
            rom[33670] = 8'h0a ;
            rom[33671] = 8'hdd ;
            rom[33672] = 8'hf3 ;
            rom[33673] = 8'hfa ;
            rom[33674] = 8'h10 ;
            rom[33675] = 8'he6 ;
            rom[33676] = 8'hf4 ;
            rom[33677] = 8'hfb ;
            rom[33678] = 8'h04 ;
            rom[33679] = 8'he4 ;
            rom[33680] = 8'hf7 ;
            rom[33681] = 8'hed ;
            rom[33682] = 8'he7 ;
            rom[33683] = 8'hdf ;
            rom[33684] = 8'h00 ;
            rom[33685] = 8'heb ;
            rom[33686] = 8'h03 ;
            rom[33687] = 8'hba ;
            rom[33688] = 8'h18 ;
            rom[33689] = 8'hf4 ;
            rom[33690] = 8'hee ;
            rom[33691] = 8'hff ;
            rom[33692] = 8'h0a ;
            rom[33693] = 8'hf0 ;
            rom[33694] = 8'hfe ;
            rom[33695] = 8'he4 ;
            rom[33696] = 8'heb ;
            rom[33697] = 8'hfe ;
            rom[33698] = 8'hdb ;
            rom[33699] = 8'hf3 ;
            rom[33700] = 8'h08 ;
            rom[33701] = 8'he8 ;
            rom[33702] = 8'hf5 ;
            rom[33703] = 8'hf9 ;
            rom[33704] = 8'hf9 ;
            rom[33705] = 8'h12 ;
            rom[33706] = 8'hfc ;
            rom[33707] = 8'hd4 ;
            rom[33708] = 8'h09 ;
            rom[33709] = 8'h08 ;
            rom[33710] = 8'hb3 ;
            rom[33711] = 8'hfa ;
            rom[33712] = 8'h14 ;
            rom[33713] = 8'hf8 ;
            rom[33714] = 8'h01 ;
            rom[33715] = 8'h09 ;
            rom[33716] = 8'h04 ;
            rom[33717] = 8'h09 ;
            rom[33718] = 8'h0a ;
            rom[33719] = 8'he8 ;
            rom[33720] = 8'h23 ;
            rom[33721] = 8'he5 ;
            rom[33722] = 8'hcf ;
            rom[33723] = 8'h1a ;
            rom[33724] = 8'h19 ;
            rom[33725] = 8'h1a ;
            rom[33726] = 8'he2 ;
            rom[33727] = 8'hd2 ;
            rom[33728] = 8'hee ;
            rom[33729] = 8'h16 ;
            rom[33730] = 8'hef ;
            rom[33731] = 8'hdf ;
            rom[33732] = 8'he6 ;
            rom[33733] = 8'he4 ;
            rom[33734] = 8'hf5 ;
            rom[33735] = 8'hfc ;
            rom[33736] = 8'hda ;
            rom[33737] = 8'h04 ;
            rom[33738] = 8'hf1 ;
            rom[33739] = 8'h0a ;
            rom[33740] = 8'hd3 ;
            rom[33741] = 8'h05 ;
            rom[33742] = 8'hc9 ;
            rom[33743] = 8'hfa ;
            rom[33744] = 8'hf0 ;
            rom[33745] = 8'hc2 ;
            rom[33746] = 8'he4 ;
            rom[33747] = 8'hb9 ;
            rom[33748] = 8'hfc ;
            rom[33749] = 8'hf0 ;
            rom[33750] = 8'h00 ;
            rom[33751] = 8'hfe ;
            rom[33752] = 8'hfe ;
            rom[33753] = 8'h0d ;
            rom[33754] = 8'hfe ;
            rom[33755] = 8'h10 ;
            rom[33756] = 8'hf3 ;
            rom[33757] = 8'hc5 ;
            rom[33758] = 8'hc2 ;
            rom[33759] = 8'he4 ;
            rom[33760] = 8'hda ;
            rom[33761] = 8'h2c ;
            rom[33762] = 8'he9 ;
            rom[33763] = 8'hf3 ;
            rom[33764] = 8'h16 ;
            rom[33765] = 8'hdd ;
            rom[33766] = 8'hf0 ;
            rom[33767] = 8'hd2 ;
            rom[33768] = 8'hf3 ;
            rom[33769] = 8'hf2 ;
            rom[33770] = 8'he4 ;
            rom[33771] = 8'hfc ;
            rom[33772] = 8'h11 ;
            rom[33773] = 8'hfc ;
            rom[33774] = 8'he1 ;
            rom[33775] = 8'hfe ;
            rom[33776] = 8'h16 ;
            rom[33777] = 8'h0a ;
            rom[33778] = 8'he9 ;
            rom[33779] = 8'h02 ;
            rom[33780] = 8'he9 ;
            rom[33781] = 8'h23 ;
            rom[33782] = 8'h15 ;
            rom[33783] = 8'h05 ;
            rom[33784] = 8'h07 ;
            rom[33785] = 8'h0b ;
            rom[33786] = 8'hec ;
            rom[33787] = 8'hef ;
            rom[33788] = 8'hdf ;
            rom[33789] = 8'h0e ;
            rom[33790] = 8'h03 ;
            rom[33791] = 8'hed ;
            rom[33792] = 8'h12 ;
            rom[33793] = 8'hfa ;
            rom[33794] = 8'h13 ;
            rom[33795] = 8'hfd ;
            rom[33796] = 8'h0c ;
            rom[33797] = 8'hed ;
            rom[33798] = 8'he3 ;
            rom[33799] = 8'hd5 ;
            rom[33800] = 8'h1e ;
            rom[33801] = 8'he6 ;
            rom[33802] = 8'h1c ;
            rom[33803] = 8'hfb ;
            rom[33804] = 8'hcf ;
            rom[33805] = 8'h11 ;
            rom[33806] = 8'hf7 ;
            rom[33807] = 8'hfe ;
            rom[33808] = 8'hdf ;
            rom[33809] = 8'hf9 ;
            rom[33810] = 8'h15 ;
            rom[33811] = 8'h04 ;
            rom[33812] = 8'he0 ;
            rom[33813] = 8'he3 ;
            rom[33814] = 8'hea ;
            rom[33815] = 8'hea ;
            rom[33816] = 8'hdb ;
            rom[33817] = 8'hfd ;
            rom[33818] = 8'hfd ;
            rom[33819] = 8'he6 ;
            rom[33820] = 8'h11 ;
            rom[33821] = 8'h0b ;
            rom[33822] = 8'h15 ;
            rom[33823] = 8'hf9 ;
            rom[33824] = 8'hf8 ;
            rom[33825] = 8'h06 ;
            rom[33826] = 8'hf6 ;
            rom[33827] = 8'h0a ;
            rom[33828] = 8'hcc ;
            rom[33829] = 8'h0b ;
            rom[33830] = 8'h00 ;
            rom[33831] = 8'h10 ;
            rom[33832] = 8'h05 ;
            rom[33833] = 8'h13 ;
            rom[33834] = 8'h04 ;
            rom[33835] = 8'h0c ;
            rom[33836] = 8'hf4 ;
            rom[33837] = 8'h14 ;
            rom[33838] = 8'he6 ;
            rom[33839] = 8'hf0 ;
            rom[33840] = 8'hc8 ;
            rom[33841] = 8'hf9 ;
            rom[33842] = 8'hf6 ;
            rom[33843] = 8'heb ;
            rom[33844] = 8'he9 ;
            rom[33845] = 8'hf4 ;
            rom[33846] = 8'hcc ;
            rom[33847] = 8'hf8 ;
            rom[33848] = 8'he3 ;
            rom[33849] = 8'hea ;
            rom[33850] = 8'hea ;
            rom[33851] = 8'hec ;
            rom[33852] = 8'h0d ;
            rom[33853] = 8'hf8 ;
            rom[33854] = 8'h0d ;
            rom[33855] = 8'hdf ;
            rom[33856] = 8'hf8 ;
            rom[33857] = 8'hec ;
            rom[33858] = 8'h00 ;
            rom[33859] = 8'hf9 ;
            rom[33860] = 8'hfb ;
            rom[33861] = 8'h2e ;
            rom[33862] = 8'hd2 ;
            rom[33863] = 8'h05 ;
            rom[33864] = 8'hff ;
            rom[33865] = 8'h0c ;
            rom[33866] = 8'hf4 ;
            rom[33867] = 8'h04 ;
            rom[33868] = 8'hf3 ;
            rom[33869] = 8'h13 ;
            rom[33870] = 8'hfe ;
            rom[33871] = 8'he8 ;
            rom[33872] = 8'hff ;
            rom[33873] = 8'hf7 ;
            rom[33874] = 8'hfc ;
            rom[33875] = 8'he5 ;
            rom[33876] = 8'h1b ;
            rom[33877] = 8'hc4 ;
            rom[33878] = 8'h10 ;
            rom[33879] = 8'h21 ;
            rom[33880] = 8'hd7 ;
            rom[33881] = 8'he7 ;
            rom[33882] = 8'hd4 ;
            rom[33883] = 8'hdd ;
            rom[33884] = 8'hc5 ;
            rom[33885] = 8'he4 ;
            rom[33886] = 8'hed ;
            rom[33887] = 8'h01 ;
            rom[33888] = 8'hee ;
            rom[33889] = 8'hfc ;
            rom[33890] = 8'hed ;
            rom[33891] = 8'hf5 ;
            rom[33892] = 8'hfc ;
            rom[33893] = 8'hf1 ;
            rom[33894] = 8'hff ;
            rom[33895] = 8'hc0 ;
            rom[33896] = 8'h09 ;
            rom[33897] = 8'h1a ;
            rom[33898] = 8'hdd ;
            rom[33899] = 8'hf2 ;
            rom[33900] = 8'he2 ;
            rom[33901] = 8'hc4 ;
            rom[33902] = 8'hfe ;
            rom[33903] = 8'hed ;
            rom[33904] = 8'hb9 ;
            rom[33905] = 8'hef ;
            rom[33906] = 8'h21 ;
            rom[33907] = 8'h12 ;
            rom[33908] = 8'hfc ;
            rom[33909] = 8'hf5 ;
            rom[33910] = 8'he6 ;
            rom[33911] = 8'hd0 ;
            rom[33912] = 8'hfa ;
            rom[33913] = 8'hdc ;
            rom[33914] = 8'hd2 ;
            rom[33915] = 8'h0a ;
            rom[33916] = 8'h14 ;
            rom[33917] = 8'he8 ;
            rom[33918] = 8'h09 ;
            rom[33919] = 8'hac ;
            rom[33920] = 8'hda ;
            rom[33921] = 8'hf5 ;
            rom[33922] = 8'hfc ;
            rom[33923] = 8'h05 ;
            rom[33924] = 8'hfd ;
            rom[33925] = 8'hf1 ;
            rom[33926] = 8'h0c ;
            rom[33927] = 8'hf4 ;
            rom[33928] = 8'hf5 ;
            rom[33929] = 8'hff ;
            rom[33930] = 8'h0e ;
            rom[33931] = 8'h1b ;
            rom[33932] = 8'hf5 ;
            rom[33933] = 8'h0a ;
            rom[33934] = 8'h1d ;
            rom[33935] = 8'hea ;
            rom[33936] = 8'h2c ;
            rom[33937] = 8'hf6 ;
            rom[33938] = 8'hff ;
            rom[33939] = 8'h1a ;
            rom[33940] = 8'h07 ;
            rom[33941] = 8'h02 ;
            rom[33942] = 8'hea ;
            rom[33943] = 8'hef ;
            rom[33944] = 8'he4 ;
            rom[33945] = 8'hce ;
            rom[33946] = 8'h0d ;
            rom[33947] = 8'hfb ;
            rom[33948] = 8'hf3 ;
            rom[33949] = 8'hdc ;
            rom[33950] = 8'hd8 ;
            rom[33951] = 8'h11 ;
            rom[33952] = 8'he7 ;
            rom[33953] = 8'h12 ;
            rom[33954] = 8'h20 ;
            rom[33955] = 8'hcb ;
            rom[33956] = 8'hed ;
            rom[33957] = 8'h08 ;
            rom[33958] = 8'hee ;
            rom[33959] = 8'hc5 ;
            rom[33960] = 8'h12 ;
            rom[33961] = 8'hfb ;
            rom[33962] = 8'hfe ;
            rom[33963] = 8'hf6 ;
            rom[33964] = 8'h04 ;
            rom[33965] = 8'h16 ;
            rom[33966] = 8'h15 ;
            rom[33967] = 8'hd3 ;
            rom[33968] = 8'he8 ;
            rom[33969] = 8'hcd ;
            rom[33970] = 8'hf9 ;
            rom[33971] = 8'he2 ;
            rom[33972] = 8'heb ;
            rom[33973] = 8'hdc ;
            rom[33974] = 8'hfd ;
            rom[33975] = 8'hef ;
            rom[33976] = 8'h00 ;
            rom[33977] = 8'hfd ;
            rom[33978] = 8'hf8 ;
            rom[33979] = 8'h07 ;
            rom[33980] = 8'h03 ;
            rom[33981] = 8'he8 ;
            rom[33982] = 8'h08 ;
            rom[33983] = 8'h10 ;
            rom[33984] = 8'h04 ;
            rom[33985] = 8'hee ;
            rom[33986] = 8'hea ;
            rom[33987] = 8'hee ;
            rom[33988] = 8'hdd ;
            rom[33989] = 8'hf9 ;
            rom[33990] = 8'hd8 ;
            rom[33991] = 8'he9 ;
            rom[33992] = 8'hf6 ;
            rom[33993] = 8'h15 ;
            rom[33994] = 8'hf4 ;
            rom[33995] = 8'h1d ;
            rom[33996] = 8'he0 ;
            rom[33997] = 8'h10 ;
            rom[33998] = 8'he9 ;
            rom[33999] = 8'h0d ;
            rom[34000] = 8'hcf ;
            rom[34001] = 8'h17 ;
            rom[34002] = 8'hfd ;
            rom[34003] = 8'h13 ;
            rom[34004] = 8'h14 ;
            rom[34005] = 8'hf4 ;
            rom[34006] = 8'hed ;
            rom[34007] = 8'hd8 ;
            rom[34008] = 8'h27 ;
            rom[34009] = 8'hed ;
            rom[34010] = 8'h13 ;
            rom[34011] = 8'h28 ;
            rom[34012] = 8'he4 ;
            rom[34013] = 8'h03 ;
            rom[34014] = 8'hf5 ;
            rom[34015] = 8'h1d ;
            rom[34016] = 8'h0c ;
            rom[34017] = 8'hfb ;
            rom[34018] = 8'h09 ;
            rom[34019] = 8'hff ;
            rom[34020] = 8'h13 ;
            rom[34021] = 8'hd8 ;
            rom[34022] = 8'hf8 ;
            rom[34023] = 8'heb ;
            rom[34024] = 8'h0c ;
            rom[34025] = 8'hec ;
            rom[34026] = 8'h03 ;
            rom[34027] = 8'h01 ;
            rom[34028] = 8'hfc ;
            rom[34029] = 8'hfe ;
            rom[34030] = 8'h13 ;
            rom[34031] = 8'hf5 ;
            rom[34032] = 8'h0e ;
            rom[34033] = 8'he3 ;
            rom[34034] = 8'h2d ;
            rom[34035] = 8'he5 ;
            rom[34036] = 8'h09 ;
            rom[34037] = 8'hf6 ;
            rom[34038] = 8'hf5 ;
            rom[34039] = 8'hed ;
            rom[34040] = 8'h10 ;
            rom[34041] = 8'h05 ;
            rom[34042] = 8'h13 ;
            rom[34043] = 8'h11 ;
            rom[34044] = 8'he4 ;
            rom[34045] = 8'hf0 ;
            rom[34046] = 8'h03 ;
            rom[34047] = 8'h03 ;
            rom[34048] = 8'h04 ;
            rom[34049] = 8'h0a ;
            rom[34050] = 8'h18 ;
            rom[34051] = 8'hec ;
            rom[34052] = 8'hda ;
            rom[34053] = 8'hfb ;
            rom[34054] = 8'h1a ;
            rom[34055] = 8'hf6 ;
            rom[34056] = 8'he8 ;
            rom[34057] = 8'h24 ;
            rom[34058] = 8'h1b ;
            rom[34059] = 8'h1e ;
            rom[34060] = 8'hf9 ;
            rom[34061] = 8'he6 ;
            rom[34062] = 8'h05 ;
            rom[34063] = 8'h01 ;
            rom[34064] = 8'hc7 ;
            rom[34065] = 8'h18 ;
            rom[34066] = 8'h0c ;
            rom[34067] = 8'h1b ;
            rom[34068] = 8'hfb ;
            rom[34069] = 8'h13 ;
            rom[34070] = 8'h34 ;
            rom[34071] = 8'h00 ;
            rom[34072] = 8'heb ;
            rom[34073] = 8'hf5 ;
            rom[34074] = 8'h00 ;
            rom[34075] = 8'h03 ;
            rom[34076] = 8'hf3 ;
            rom[34077] = 8'hf5 ;
            rom[34078] = 8'hfc ;
            rom[34079] = 8'hf8 ;
            rom[34080] = 8'h06 ;
            rom[34081] = 8'hfb ;
            rom[34082] = 8'hde ;
            rom[34083] = 8'h17 ;
            rom[34084] = 8'h1b ;
            rom[34085] = 8'hec ;
            rom[34086] = 8'hee ;
            rom[34087] = 8'hee ;
            rom[34088] = 8'hf9 ;
            rom[34089] = 8'he9 ;
            rom[34090] = 8'h02 ;
            rom[34091] = 8'h03 ;
            rom[34092] = 8'he6 ;
            rom[34093] = 8'hf4 ;
            rom[34094] = 8'hff ;
            rom[34095] = 8'hd0 ;
            rom[34096] = 8'hea ;
            rom[34097] = 8'hef ;
            rom[34098] = 8'hf4 ;
            rom[34099] = 8'hf2 ;
            rom[34100] = 8'hc6 ;
            rom[34101] = 8'h0f ;
            rom[34102] = 8'hff ;
            rom[34103] = 8'hf2 ;
            rom[34104] = 8'hef ;
            rom[34105] = 8'h1f ;
            rom[34106] = 8'he0 ;
            rom[34107] = 8'h15 ;
            rom[34108] = 8'hf9 ;
            rom[34109] = 8'hfc ;
            rom[34110] = 8'hf9 ;
            rom[34111] = 8'hf6 ;
            rom[34112] = 8'h08 ;
            rom[34113] = 8'hde ;
            rom[34114] = 8'h27 ;
            rom[34115] = 8'hd4 ;
            rom[34116] = 8'hfe ;
            rom[34117] = 8'he6 ;
            rom[34118] = 8'hcc ;
            rom[34119] = 8'hf2 ;
            rom[34120] = 8'hf6 ;
            rom[34121] = 8'h0c ;
            rom[34122] = 8'hde ;
            rom[34123] = 8'h24 ;
            rom[34124] = 8'hc0 ;
            rom[34125] = 8'h1e ;
            rom[34126] = 8'hf0 ;
            rom[34127] = 8'h0f ;
            rom[34128] = 8'h11 ;
            rom[34129] = 8'h0d ;
            rom[34130] = 8'hcc ;
            rom[34131] = 8'hed ;
            rom[34132] = 8'h07 ;
            rom[34133] = 8'hdc ;
            rom[34134] = 8'he0 ;
            rom[34135] = 8'hea ;
            rom[34136] = 8'hdd ;
            rom[34137] = 8'h0d ;
            rom[34138] = 8'he3 ;
            rom[34139] = 8'h07 ;
            rom[34140] = 8'he6 ;
            rom[34141] = 8'hfc ;
            rom[34142] = 8'he4 ;
            rom[34143] = 8'he8 ;
            rom[34144] = 8'hf7 ;
            rom[34145] = 8'h00 ;
            rom[34146] = 8'h13 ;
            rom[34147] = 8'h09 ;
            rom[34148] = 8'h1b ;
            rom[34149] = 8'he3 ;
            rom[34150] = 8'h12 ;
            rom[34151] = 8'h0c ;
            rom[34152] = 8'he2 ;
            rom[34153] = 8'h0b ;
            rom[34154] = 8'hf0 ;
            rom[34155] = 8'hf7 ;
            rom[34156] = 8'he5 ;
            rom[34157] = 8'h04 ;
            rom[34158] = 8'h0a ;
            rom[34159] = 8'h13 ;
            rom[34160] = 8'h01 ;
            rom[34161] = 8'hfb ;
            rom[34162] = 8'h0d ;
            rom[34163] = 8'hfa ;
            rom[34164] = 8'h1d ;
            rom[34165] = 8'heb ;
            rom[34166] = 8'hfd ;
            rom[34167] = 8'h11 ;
            rom[34168] = 8'hff ;
            rom[34169] = 8'h26 ;
            rom[34170] = 8'he8 ;
            rom[34171] = 8'hf6 ;
            rom[34172] = 8'h20 ;
            rom[34173] = 8'h00 ;
            rom[34174] = 8'h01 ;
            rom[34175] = 8'hf6 ;
            rom[34176] = 8'hfb ;
            rom[34177] = 8'hfc ;
            rom[34178] = 8'hfa ;
            rom[34179] = 8'hcf ;
            rom[34180] = 8'hca ;
            rom[34181] = 8'h18 ;
            rom[34182] = 8'h02 ;
            rom[34183] = 8'h09 ;
            rom[34184] = 8'hfb ;
            rom[34185] = 8'hfc ;
            rom[34186] = 8'hfb ;
            rom[34187] = 8'hd0 ;
            rom[34188] = 8'hf2 ;
            rom[34189] = 8'hf6 ;
            rom[34190] = 8'h16 ;
            rom[34191] = 8'hdc ;
            rom[34192] = 8'h0d ;
            rom[34193] = 8'h05 ;
            rom[34194] = 8'hff ;
            rom[34195] = 8'h00 ;
            rom[34196] = 8'hea ;
            rom[34197] = 8'hf5 ;
            rom[34198] = 8'he9 ;
            rom[34199] = 8'hcf ;
            rom[34200] = 8'hea ;
            rom[34201] = 8'hfc ;
            rom[34202] = 8'ha3 ;
            rom[34203] = 8'h12 ;
            rom[34204] = 8'h13 ;
            rom[34205] = 8'hdd ;
            rom[34206] = 8'hed ;
            rom[34207] = 8'he7 ;
            rom[34208] = 8'h02 ;
            rom[34209] = 8'h17 ;
            rom[34210] = 8'h04 ;
            rom[34211] = 8'hf6 ;
            rom[34212] = 8'hff ;
            rom[34213] = 8'hf7 ;
            rom[34214] = 8'h02 ;
            rom[34215] = 8'hf3 ;
            rom[34216] = 8'hb7 ;
            rom[34217] = 8'he4 ;
            rom[34218] = 8'h10 ;
            rom[34219] = 8'h06 ;
            rom[34220] = 8'he9 ;
            rom[34221] = 8'ha4 ;
            rom[34222] = 8'he9 ;
            rom[34223] = 8'hfe ;
            rom[34224] = 8'hfb ;
            rom[34225] = 8'h03 ;
            rom[34226] = 8'hb6 ;
            rom[34227] = 8'h10 ;
            rom[34228] = 8'had ;
            rom[34229] = 8'h0a ;
            rom[34230] = 8'h23 ;
            rom[34231] = 8'hf8 ;
            rom[34232] = 8'h03 ;
            rom[34233] = 8'hff ;
            rom[34234] = 8'h04 ;
            rom[34235] = 8'hf5 ;
            rom[34236] = 8'hf8 ;
            rom[34237] = 8'hec ;
            rom[34238] = 8'h18 ;
            rom[34239] = 8'hfd ;
            rom[34240] = 8'h01 ;
            rom[34241] = 8'h03 ;
            rom[34242] = 8'h05 ;
            rom[34243] = 8'hfa ;
            rom[34244] = 8'hd6 ;
            rom[34245] = 8'hfb ;
            rom[34246] = 8'h16 ;
            rom[34247] = 8'h01 ;
            rom[34248] = 8'hf7 ;
            rom[34249] = 8'hfa ;
            rom[34250] = 8'hf2 ;
            rom[34251] = 8'hd3 ;
            rom[34252] = 8'hdc ;
            rom[34253] = 8'hf0 ;
            rom[34254] = 8'he7 ;
            rom[34255] = 8'hf8 ;
            rom[34256] = 8'hf6 ;
            rom[34257] = 8'hd1 ;
            rom[34258] = 8'h08 ;
            rom[34259] = 8'hd0 ;
            rom[34260] = 8'hf4 ;
            rom[34261] = 8'he8 ;
            rom[34262] = 8'hf4 ;
            rom[34263] = 8'h0c ;
            rom[34264] = 8'h15 ;
            rom[34265] = 8'heb ;
            rom[34266] = 8'h11 ;
            rom[34267] = 8'hf0 ;
            rom[34268] = 8'hfd ;
            rom[34269] = 8'hfe ;
            rom[34270] = 8'hc2 ;
            rom[34271] = 8'he0 ;
            rom[34272] = 8'he5 ;
            rom[34273] = 8'hf7 ;
            rom[34274] = 8'hfd ;
            rom[34275] = 8'h0f ;
            rom[34276] = 8'hfc ;
            rom[34277] = 8'h08 ;
            rom[34278] = 8'h19 ;
            rom[34279] = 8'h1e ;
            rom[34280] = 8'haa ;
            rom[34281] = 8'hfd ;
            rom[34282] = 8'hff ;
            rom[34283] = 8'hfc ;
            rom[34284] = 8'h0f ;
            rom[34285] = 8'hfb ;
            rom[34286] = 8'hf5 ;
            rom[34287] = 8'h13 ;
            rom[34288] = 8'h15 ;
            rom[34289] = 8'hd4 ;
            rom[34290] = 8'h0f ;
            rom[34291] = 8'he6 ;
            rom[34292] = 8'hf4 ;
            rom[34293] = 8'hfc ;
            rom[34294] = 8'hfc ;
            rom[34295] = 8'h0a ;
            rom[34296] = 8'hfa ;
            rom[34297] = 8'hf0 ;
            rom[34298] = 8'h02 ;
            rom[34299] = 8'hff ;
            rom[34300] = 8'hc9 ;
            rom[34301] = 8'hf0 ;
            rom[34302] = 8'h01 ;
            rom[34303] = 8'h23 ;
            rom[34304] = 8'hda ;
            rom[34305] = 8'hf0 ;
            rom[34306] = 8'h1c ;
            rom[34307] = 8'hff ;
            rom[34308] = 8'hb2 ;
            rom[34309] = 8'h26 ;
            rom[34310] = 8'hfb ;
            rom[34311] = 8'h0a ;
            rom[34312] = 8'h27 ;
            rom[34313] = 8'h04 ;
            rom[34314] = 8'hd9 ;
            rom[34315] = 8'h0b ;
            rom[34316] = 8'h15 ;
            rom[34317] = 8'hde ;
            rom[34318] = 8'hfb ;
            rom[34319] = 8'h17 ;
            rom[34320] = 8'he7 ;
            rom[34321] = 8'h21 ;
            rom[34322] = 8'hf5 ;
            rom[34323] = 8'h1c ;
            rom[34324] = 8'h1b ;
            rom[34325] = 8'hdc ;
            rom[34326] = 8'h02 ;
            rom[34327] = 8'hf9 ;
            rom[34328] = 8'hf1 ;
            rom[34329] = 8'h02 ;
            rom[34330] = 8'hf9 ;
            rom[34331] = 8'hfd ;
            rom[34332] = 8'h01 ;
            rom[34333] = 8'h00 ;
            rom[34334] = 8'hf6 ;
            rom[34335] = 8'hf7 ;
            rom[34336] = 8'hfb ;
            rom[34337] = 8'he6 ;
            rom[34338] = 8'hed ;
            rom[34339] = 8'hfd ;
            rom[34340] = 8'h2b ;
            rom[34341] = 8'he5 ;
            rom[34342] = 8'h01 ;
            rom[34343] = 8'he5 ;
            rom[34344] = 8'hf5 ;
            rom[34345] = 8'hce ;
            rom[34346] = 8'hfc ;
            rom[34347] = 8'h0b ;
            rom[34348] = 8'he6 ;
            rom[34349] = 8'hee ;
            rom[34350] = 8'hda ;
            rom[34351] = 8'hf7 ;
            rom[34352] = 8'h0d ;
            rom[34353] = 8'h0c ;
            rom[34354] = 8'hfd ;
            rom[34355] = 8'h0c ;
            rom[34356] = 8'hf3 ;
            rom[34357] = 8'h0a ;
            rom[34358] = 8'h17 ;
            rom[34359] = 8'hd4 ;
            rom[34360] = 8'h0b ;
            rom[34361] = 8'h11 ;
            rom[34362] = 8'hc0 ;
            rom[34363] = 8'h03 ;
            rom[34364] = 8'hf2 ;
            rom[34365] = 8'hf5 ;
            rom[34366] = 8'h11 ;
            rom[34367] = 8'hec ;
            rom[34368] = 8'h1b ;
            rom[34369] = 8'h11 ;
            rom[34370] = 8'h01 ;
            rom[34371] = 8'h14 ;
            rom[34372] = 8'h07 ;
            rom[34373] = 8'h04 ;
            rom[34374] = 8'h29 ;
            rom[34375] = 8'hff ;
            rom[34376] = 8'he7 ;
            rom[34377] = 8'hfb ;
            rom[34378] = 8'hec ;
            rom[34379] = 8'h16 ;
            rom[34380] = 8'hd3 ;
            rom[34381] = 8'hed ;
            rom[34382] = 8'hf1 ;
            rom[34383] = 8'h01 ;
            rom[34384] = 8'h21 ;
            rom[34385] = 8'h14 ;
            rom[34386] = 8'h0a ;
            rom[34387] = 8'he3 ;
            rom[34388] = 8'h05 ;
            rom[34389] = 8'h04 ;
            rom[34390] = 8'h15 ;
            rom[34391] = 8'heb ;
            rom[34392] = 8'hf9 ;
            rom[34393] = 8'hfa ;
            rom[34394] = 8'hc2 ;
            rom[34395] = 8'hed ;
            rom[34396] = 8'h12 ;
            rom[34397] = 8'he2 ;
            rom[34398] = 8'h0d ;
            rom[34399] = 8'hcf ;
            rom[34400] = 8'hee ;
            rom[34401] = 8'hf7 ;
            rom[34402] = 8'hc3 ;
            rom[34403] = 8'h12 ;
            rom[34404] = 8'hf5 ;
            rom[34405] = 8'hfb ;
            rom[34406] = 8'hf4 ;
            rom[34407] = 8'h10 ;
            rom[34408] = 8'h0c ;
            rom[34409] = 8'h08 ;
            rom[34410] = 8'h1b ;
            rom[34411] = 8'hf4 ;
            rom[34412] = 8'hf6 ;
            rom[34413] = 8'hf4 ;
            rom[34414] = 8'hf0 ;
            rom[34415] = 8'hed ;
            rom[34416] = 8'h14 ;
            rom[34417] = 8'hfe ;
            rom[34418] = 8'hf6 ;
            rom[34419] = 8'hfa ;
            rom[34420] = 8'he8 ;
            rom[34421] = 8'he4 ;
            rom[34422] = 8'h02 ;
            rom[34423] = 8'h17 ;
            rom[34424] = 8'hef ;
            rom[34425] = 8'he2 ;
            rom[34426] = 8'hda ;
            rom[34427] = 8'hff ;
            rom[34428] = 8'hf6 ;
            rom[34429] = 8'hff ;
            rom[34430] = 8'hd8 ;
            rom[34431] = 8'h15 ;
            rom[34432] = 8'hf4 ;
            rom[34433] = 8'h13 ;
            rom[34434] = 8'he1 ;
            rom[34435] = 8'h26 ;
            rom[34436] = 8'h04 ;
            rom[34437] = 8'h07 ;
            rom[34438] = 8'h21 ;
            rom[34439] = 8'hec ;
            rom[34440] = 8'h00 ;
            rom[34441] = 8'hf0 ;
            rom[34442] = 8'he9 ;
            rom[34443] = 8'h11 ;
            rom[34444] = 8'hfb ;
            rom[34445] = 8'hce ;
            rom[34446] = 8'h14 ;
            rom[34447] = 8'h00 ;
            rom[34448] = 8'he7 ;
            rom[34449] = 8'h13 ;
            rom[34450] = 8'he5 ;
            rom[34451] = 8'h0d ;
            rom[34452] = 8'h03 ;
            rom[34453] = 8'h03 ;
            rom[34454] = 8'h13 ;
            rom[34455] = 8'h14 ;
            rom[34456] = 8'h11 ;
            rom[34457] = 8'hea ;
            rom[34458] = 8'hfa ;
            rom[34459] = 8'hf0 ;
            rom[34460] = 8'h0a ;
            rom[34461] = 8'h07 ;
            rom[34462] = 8'h11 ;
            rom[34463] = 8'h12 ;
            rom[34464] = 8'hed ;
            rom[34465] = 8'hfe ;
            rom[34466] = 8'hca ;
            rom[34467] = 8'hee ;
            rom[34468] = 8'hfb ;
            rom[34469] = 8'h03 ;
            rom[34470] = 8'hd4 ;
            rom[34471] = 8'h09 ;
            rom[34472] = 8'he5 ;
            rom[34473] = 8'hf8 ;
            rom[34474] = 8'h13 ;
            rom[34475] = 8'h1e ;
            rom[34476] = 8'h0e ;
            rom[34477] = 8'hce ;
            rom[34478] = 8'hef ;
            rom[34479] = 8'hf7 ;
            rom[34480] = 8'hff ;
            rom[34481] = 8'h10 ;
            rom[34482] = 8'h01 ;
            rom[34483] = 8'hf0 ;
            rom[34484] = 8'hc2 ;
            rom[34485] = 8'hf9 ;
            rom[34486] = 8'hf8 ;
            rom[34487] = 8'hf0 ;
            rom[34488] = 8'hf2 ;
            rom[34489] = 8'h0b ;
            rom[34490] = 8'hf6 ;
            rom[34491] = 8'hff ;
            rom[34492] = 8'h16 ;
            rom[34493] = 8'h0e ;
            rom[34494] = 8'h1e ;
            rom[34495] = 8'hfe ;
            rom[34496] = 8'hd4 ;
            rom[34497] = 8'he9 ;
            rom[34498] = 8'h07 ;
            rom[34499] = 8'he3 ;
            rom[34500] = 8'hdf ;
            rom[34501] = 8'hf7 ;
            rom[34502] = 8'hd4 ;
            rom[34503] = 8'h00 ;
            rom[34504] = 8'h06 ;
            rom[34505] = 8'h08 ;
            rom[34506] = 8'hfb ;
            rom[34507] = 8'hf0 ;
            rom[34508] = 8'h03 ;
            rom[34509] = 8'hee ;
            rom[34510] = 8'hf3 ;
            rom[34511] = 8'hd7 ;
            rom[34512] = 8'heb ;
            rom[34513] = 8'h08 ;
            rom[34514] = 8'h04 ;
            rom[34515] = 8'hf8 ;
            rom[34516] = 8'h0b ;
            rom[34517] = 8'hdc ;
            rom[34518] = 8'h09 ;
            rom[34519] = 8'he2 ;
            rom[34520] = 8'h02 ;
            rom[34521] = 8'h1d ;
            rom[34522] = 8'h1e ;
            rom[34523] = 8'h05 ;
            rom[34524] = 8'h0c ;
            rom[34525] = 8'h04 ;
            rom[34526] = 8'h15 ;
            rom[34527] = 8'hd3 ;
            rom[34528] = 8'hef ;
            rom[34529] = 8'h13 ;
            rom[34530] = 8'hfc ;
            rom[34531] = 8'hf3 ;
            rom[34532] = 8'h00 ;
            rom[34533] = 8'he7 ;
            rom[34534] = 8'hf7 ;
            rom[34535] = 8'hfd ;
            rom[34536] = 8'hf7 ;
            rom[34537] = 8'h25 ;
            rom[34538] = 8'hbb ;
            rom[34539] = 8'h03 ;
            rom[34540] = 8'h11 ;
            rom[34541] = 8'hfb ;
            rom[34542] = 8'he0 ;
            rom[34543] = 8'h24 ;
            rom[34544] = 8'h05 ;
            rom[34545] = 8'hf8 ;
            rom[34546] = 8'hed ;
            rom[34547] = 8'hf9 ;
            rom[34548] = 8'h09 ;
            rom[34549] = 8'h0e ;
            rom[34550] = 8'h23 ;
            rom[34551] = 8'h19 ;
            rom[34552] = 8'h0a ;
            rom[34553] = 8'hfa ;
            rom[34554] = 8'hed ;
            rom[34555] = 8'h26 ;
            rom[34556] = 8'hf6 ;
            rom[34557] = 8'h10 ;
            rom[34558] = 8'hfb ;
            rom[34559] = 8'h02 ;
            rom[34560] = 8'h1e ;
            rom[34561] = 8'hf1 ;
            rom[34562] = 8'h0d ;
            rom[34563] = 8'h0f ;
            rom[34564] = 8'h07 ;
            rom[34565] = 8'hf9 ;
            rom[34566] = 8'h02 ;
            rom[34567] = 8'hdf ;
            rom[34568] = 8'h05 ;
            rom[34569] = 8'hec ;
            rom[34570] = 8'hee ;
            rom[34571] = 8'hf7 ;
            rom[34572] = 8'h06 ;
            rom[34573] = 8'hda ;
            rom[34574] = 8'h15 ;
            rom[34575] = 8'hee ;
            rom[34576] = 8'h14 ;
            rom[34577] = 8'heb ;
            rom[34578] = 8'hfc ;
            rom[34579] = 8'h15 ;
            rom[34580] = 8'hd6 ;
            rom[34581] = 8'hc7 ;
            rom[34582] = 8'h06 ;
            rom[34583] = 8'h0d ;
            rom[34584] = 8'hec ;
            rom[34585] = 8'h1a ;
            rom[34586] = 8'hf2 ;
            rom[34587] = 8'hee ;
            rom[34588] = 8'he3 ;
            rom[34589] = 8'h01 ;
            rom[34590] = 8'h0d ;
            rom[34591] = 8'hd1 ;
            rom[34592] = 8'h0a ;
            rom[34593] = 8'h0a ;
            rom[34594] = 8'hf8 ;
            rom[34595] = 8'hf2 ;
            rom[34596] = 8'hf4 ;
            rom[34597] = 8'h38 ;
            rom[34598] = 8'h01 ;
            rom[34599] = 8'h1a ;
            rom[34600] = 8'hd9 ;
            rom[34601] = 8'hc9 ;
            rom[34602] = 8'h2a ;
            rom[34603] = 8'h0c ;
            rom[34604] = 8'h0e ;
            rom[34605] = 8'h06 ;
            rom[34606] = 8'h0b ;
            rom[34607] = 8'h04 ;
            rom[34608] = 8'he7 ;
            rom[34609] = 8'h21 ;
            rom[34610] = 8'h07 ;
            rom[34611] = 8'h03 ;
            rom[34612] = 8'h0b ;
            rom[34613] = 8'hee ;
            rom[34614] = 8'hf7 ;
            rom[34615] = 8'he5 ;
            rom[34616] = 8'hf6 ;
            rom[34617] = 8'h2c ;
            rom[34618] = 8'h17 ;
            rom[34619] = 8'hbe ;
            rom[34620] = 8'hde ;
            rom[34621] = 8'h00 ;
            rom[34622] = 8'hf7 ;
            rom[34623] = 8'h16 ;
            rom[34624] = 8'hd6 ;
            rom[34625] = 8'he3 ;
            rom[34626] = 8'h19 ;
            rom[34627] = 8'hf0 ;
            rom[34628] = 8'he2 ;
            rom[34629] = 8'h02 ;
            rom[34630] = 8'he1 ;
            rom[34631] = 8'he8 ;
            rom[34632] = 8'h02 ;
            rom[34633] = 8'hef ;
            rom[34634] = 8'hfc ;
            rom[34635] = 8'hdb ;
            rom[34636] = 8'hea ;
            rom[34637] = 8'heb ;
            rom[34638] = 8'hf1 ;
            rom[34639] = 8'he6 ;
            rom[34640] = 8'h1f ;
            rom[34641] = 8'hd8 ;
            rom[34642] = 8'h12 ;
            rom[34643] = 8'hfe ;
            rom[34644] = 8'hf0 ;
            rom[34645] = 8'h01 ;
            rom[34646] = 8'h09 ;
            rom[34647] = 8'h17 ;
            rom[34648] = 8'h0b ;
            rom[34649] = 8'h0d ;
            rom[34650] = 8'h13 ;
            rom[34651] = 8'h10 ;
            rom[34652] = 8'hfb ;
            rom[34653] = 8'hed ;
            rom[34654] = 8'h03 ;
            rom[34655] = 8'hea ;
            rom[34656] = 8'h00 ;
            rom[34657] = 8'hf4 ;
            rom[34658] = 8'hfe ;
            rom[34659] = 8'h29 ;
            rom[34660] = 8'hf3 ;
            rom[34661] = 8'h0c ;
            rom[34662] = 8'hf1 ;
            rom[34663] = 8'hf3 ;
            rom[34664] = 8'hdf ;
            rom[34665] = 8'he3 ;
            rom[34666] = 8'hf8 ;
            rom[34667] = 8'h22 ;
            rom[34668] = 8'hf1 ;
            rom[34669] = 8'h0e ;
            rom[34670] = 8'hf3 ;
            rom[34671] = 8'hfb ;
            rom[34672] = 8'hea ;
            rom[34673] = 8'hed ;
            rom[34674] = 8'h08 ;
            rom[34675] = 8'hfb ;
            rom[34676] = 8'h03 ;
            rom[34677] = 8'h1b ;
            rom[34678] = 8'hf9 ;
            rom[34679] = 8'h12 ;
            rom[34680] = 8'h24 ;
            rom[34681] = 8'hfd ;
            rom[34682] = 8'h0e ;
            rom[34683] = 8'h01 ;
            rom[34684] = 8'h00 ;
            rom[34685] = 8'hf8 ;
            rom[34686] = 8'hfb ;
            rom[34687] = 8'h04 ;
            rom[34688] = 8'hed ;
            rom[34689] = 8'hf1 ;
            rom[34690] = 8'h0c ;
            rom[34691] = 8'h08 ;
            rom[34692] = 8'hf2 ;
            rom[34693] = 8'h0a ;
            rom[34694] = 8'h19 ;
            rom[34695] = 8'heb ;
            rom[34696] = 8'h19 ;
            rom[34697] = 8'hf9 ;
            rom[34698] = 8'hf0 ;
            rom[34699] = 8'h00 ;
            rom[34700] = 8'h11 ;
            rom[34701] = 8'hec ;
            rom[34702] = 8'h0a ;
            rom[34703] = 8'he5 ;
            rom[34704] = 8'h02 ;
            rom[34705] = 8'hc6 ;
            rom[34706] = 8'hf7 ;
            rom[34707] = 8'hc3 ;
            rom[34708] = 8'h0f ;
            rom[34709] = 8'h05 ;
            rom[34710] = 8'hf6 ;
            rom[34711] = 8'he7 ;
            rom[34712] = 8'h08 ;
            rom[34713] = 8'h02 ;
            rom[34714] = 8'h09 ;
            rom[34715] = 8'hf6 ;
            rom[34716] = 8'h02 ;
            rom[34717] = 8'hf4 ;
            rom[34718] = 8'h1b ;
            rom[34719] = 8'h22 ;
            rom[34720] = 8'h1c ;
            rom[34721] = 8'hd4 ;
            rom[34722] = 8'hd3 ;
            rom[34723] = 8'h1f ;
            rom[34724] = 8'hfd ;
            rom[34725] = 8'h04 ;
            rom[34726] = 8'h1b ;
            rom[34727] = 8'h12 ;
            rom[34728] = 8'h0f ;
            rom[34729] = 8'hee ;
            rom[34730] = 8'h1a ;
            rom[34731] = 8'hf4 ;
            rom[34732] = 8'h0c ;
            rom[34733] = 8'hf0 ;
            rom[34734] = 8'hfc ;
            rom[34735] = 8'hef ;
            rom[34736] = 8'hf0 ;
            rom[34737] = 8'h13 ;
            rom[34738] = 8'h0c ;
            rom[34739] = 8'h26 ;
            rom[34740] = 8'hf1 ;
            rom[34741] = 8'h13 ;
            rom[34742] = 8'h0b ;
            rom[34743] = 8'hd8 ;
            rom[34744] = 8'h12 ;
            rom[34745] = 8'hfc ;
            rom[34746] = 8'hff ;
            rom[34747] = 8'h11 ;
            rom[34748] = 8'h01 ;
            rom[34749] = 8'h28 ;
            rom[34750] = 8'hdb ;
            rom[34751] = 8'hf5 ;
            rom[34752] = 8'hfc ;
            rom[34753] = 8'h24 ;
            rom[34754] = 8'he6 ;
            rom[34755] = 8'hdd ;
            rom[34756] = 8'h14 ;
            rom[34757] = 8'heb ;
            rom[34758] = 8'hf8 ;
            rom[34759] = 8'h18 ;
            rom[34760] = 8'hf4 ;
            rom[34761] = 8'h00 ;
            rom[34762] = 8'h1a ;
            rom[34763] = 8'hfb ;
            rom[34764] = 8'hfd ;
            rom[34765] = 8'hd0 ;
            rom[34766] = 8'hd0 ;
            rom[34767] = 8'hd5 ;
            rom[34768] = 8'h20 ;
            rom[34769] = 8'hd2 ;
            rom[34770] = 8'h18 ;
            rom[34771] = 8'h0e ;
            rom[34772] = 8'hd7 ;
            rom[34773] = 8'hef ;
            rom[34774] = 8'h23 ;
            rom[34775] = 8'hcf ;
            rom[34776] = 8'h1e ;
            rom[34777] = 8'h0b ;
            rom[34778] = 8'h1f ;
            rom[34779] = 8'h11 ;
            rom[34780] = 8'h00 ;
            rom[34781] = 8'hf3 ;
            rom[34782] = 8'he9 ;
            rom[34783] = 8'hf2 ;
            rom[34784] = 8'hd9 ;
            rom[34785] = 8'h33 ;
            rom[34786] = 8'hfb ;
            rom[34787] = 8'hdc ;
            rom[34788] = 8'h00 ;
            rom[34789] = 8'hd5 ;
            rom[34790] = 8'he9 ;
            rom[34791] = 8'hdc ;
            rom[34792] = 8'h02 ;
            rom[34793] = 8'hec ;
            rom[34794] = 8'hfa ;
            rom[34795] = 8'h15 ;
            rom[34796] = 8'hdb ;
            rom[34797] = 8'h0c ;
            rom[34798] = 8'hd9 ;
            rom[34799] = 8'h27 ;
            rom[34800] = 8'h13 ;
            rom[34801] = 8'hff ;
            rom[34802] = 8'hf4 ;
            rom[34803] = 8'h10 ;
            rom[34804] = 8'hf6 ;
            rom[34805] = 8'h20 ;
            rom[34806] = 8'h06 ;
            rom[34807] = 8'he5 ;
            rom[34808] = 8'he7 ;
            rom[34809] = 8'h07 ;
            rom[34810] = 8'h14 ;
            rom[34811] = 8'h03 ;
            rom[34812] = 8'he4 ;
            rom[34813] = 8'hf4 ;
            rom[34814] = 8'hff ;
            rom[34815] = 8'h19 ;
            rom[34816] = 8'heb ;
            rom[34817] = 8'h0c ;
            rom[34818] = 8'hfb ;
            rom[34819] = 8'h10 ;
            rom[34820] = 8'h0e ;
            rom[34821] = 8'hf2 ;
            rom[34822] = 8'h12 ;
            rom[34823] = 8'he3 ;
            rom[34824] = 8'he9 ;
            rom[34825] = 8'h04 ;
            rom[34826] = 8'hc8 ;
            rom[34827] = 8'h11 ;
            rom[34828] = 8'hf0 ;
            rom[34829] = 8'hf5 ;
            rom[34830] = 8'hb8 ;
            rom[34831] = 8'h11 ;
            rom[34832] = 8'h17 ;
            rom[34833] = 8'h09 ;
            rom[34834] = 8'he5 ;
            rom[34835] = 8'h02 ;
            rom[34836] = 8'h12 ;
            rom[34837] = 8'h22 ;
            rom[34838] = 8'hdc ;
            rom[34839] = 8'h19 ;
            rom[34840] = 8'h0a ;
            rom[34841] = 8'h07 ;
            rom[34842] = 8'hf1 ;
            rom[34843] = 8'h08 ;
            rom[34844] = 8'he7 ;
            rom[34845] = 8'he4 ;
            rom[34846] = 8'h04 ;
            rom[34847] = 8'h18 ;
            rom[34848] = 8'h08 ;
            rom[34849] = 8'h1c ;
            rom[34850] = 8'hd6 ;
            rom[34851] = 8'hec ;
            rom[34852] = 8'hfb ;
            rom[34853] = 8'hd8 ;
            rom[34854] = 8'hfe ;
            rom[34855] = 8'h06 ;
            rom[34856] = 8'h0c ;
            rom[34857] = 8'he3 ;
            rom[34858] = 8'h0f ;
            rom[34859] = 8'h10 ;
            rom[34860] = 8'h1a ;
            rom[34861] = 8'hce ;
            rom[34862] = 8'hfc ;
            rom[34863] = 8'h05 ;
            rom[34864] = 8'h06 ;
            rom[34865] = 8'hf5 ;
            rom[34866] = 8'h1a ;
            rom[34867] = 8'hfe ;
            rom[34868] = 8'he1 ;
            rom[34869] = 8'hfd ;
            rom[34870] = 8'h11 ;
            rom[34871] = 8'h02 ;
            rom[34872] = 8'hd0 ;
            rom[34873] = 8'h12 ;
            rom[34874] = 8'h03 ;
            rom[34875] = 8'h07 ;
            rom[34876] = 8'heb ;
            rom[34877] = 8'h0c ;
            rom[34878] = 8'hf6 ;
            rom[34879] = 8'hec ;
            rom[34880] = 8'hc9 ;
            rom[34881] = 8'heb ;
            rom[34882] = 8'h11 ;
            rom[34883] = 8'he0 ;
            rom[34884] = 8'hea ;
            rom[34885] = 8'h11 ;
            rom[34886] = 8'h02 ;
            rom[34887] = 8'hf7 ;
            rom[34888] = 8'hdb ;
            rom[34889] = 8'h0b ;
            rom[34890] = 8'h0c ;
            rom[34891] = 8'hf5 ;
            rom[34892] = 8'h07 ;
            rom[34893] = 8'hcd ;
            rom[34894] = 8'hf8 ;
            rom[34895] = 8'h05 ;
            rom[34896] = 8'h07 ;
            rom[34897] = 8'h16 ;
            rom[34898] = 8'hdd ;
            rom[34899] = 8'hf1 ;
            rom[34900] = 8'hf3 ;
            rom[34901] = 8'hd1 ;
            rom[34902] = 8'h01 ;
            rom[34903] = 8'h0b ;
            rom[34904] = 8'hf0 ;
            rom[34905] = 8'h18 ;
            rom[34906] = 8'h08 ;
            rom[34907] = 8'he1 ;
            rom[34908] = 8'h07 ;
            rom[34909] = 8'h02 ;
            rom[34910] = 8'h03 ;
            rom[34911] = 8'hd5 ;
            rom[34912] = 8'h12 ;
            rom[34913] = 8'h04 ;
            rom[34914] = 8'he3 ;
            rom[34915] = 8'hf9 ;
            rom[34916] = 8'h06 ;
            rom[34917] = 8'hfe ;
            rom[34918] = 8'h08 ;
            rom[34919] = 8'he4 ;
            rom[34920] = 8'h02 ;
            rom[34921] = 8'hfa ;
            rom[34922] = 8'he5 ;
            rom[34923] = 8'h12 ;
            rom[34924] = 8'hdb ;
            rom[34925] = 8'he7 ;
            rom[34926] = 8'hdb ;
            rom[34927] = 8'h00 ;
            rom[34928] = 8'he7 ;
            rom[34929] = 8'hf4 ;
            rom[34930] = 8'h0e ;
            rom[34931] = 8'hf9 ;
            rom[34932] = 8'h0d ;
            rom[34933] = 8'h1c ;
            rom[34934] = 8'h08 ;
            rom[34935] = 8'h0a ;
            rom[34936] = 8'h13 ;
            rom[34937] = 8'h16 ;
            rom[34938] = 8'hcd ;
            rom[34939] = 8'h09 ;
            rom[34940] = 8'h0d ;
            rom[34941] = 8'h08 ;
            rom[34942] = 8'hf1 ;
            rom[34943] = 8'h01 ;
            rom[34944] = 8'h0e ;
            rom[34945] = 8'hf2 ;
            rom[34946] = 8'h10 ;
            rom[34947] = 8'hd5 ;
            rom[34948] = 8'hd1 ;
            rom[34949] = 8'hf4 ;
            rom[34950] = 8'h1e ;
            rom[34951] = 8'hf8 ;
            rom[34952] = 8'hf8 ;
            rom[34953] = 8'hdd ;
            rom[34954] = 8'hfe ;
            rom[34955] = 8'hff ;
            rom[34956] = 8'h24 ;
            rom[34957] = 8'hf2 ;
            rom[34958] = 8'hf1 ;
            rom[34959] = 8'hf5 ;
            rom[34960] = 8'h09 ;
            rom[34961] = 8'h09 ;
            rom[34962] = 8'hfe ;
            rom[34963] = 8'h06 ;
            rom[34964] = 8'hec ;
            rom[34965] = 8'hd0 ;
            rom[34966] = 8'hfb ;
            rom[34967] = 8'he3 ;
            rom[34968] = 8'hcf ;
            rom[34969] = 8'hfe ;
            rom[34970] = 8'he1 ;
            rom[34971] = 8'hed ;
            rom[34972] = 8'h09 ;
            rom[34973] = 8'hdb ;
            rom[34974] = 8'hf3 ;
            rom[34975] = 8'h0c ;
            rom[34976] = 8'hf1 ;
            rom[34977] = 8'h14 ;
            rom[34978] = 8'he9 ;
            rom[34979] = 8'hff ;
            rom[34980] = 8'h12 ;
            rom[34981] = 8'h09 ;
            rom[34982] = 8'h0f ;
            rom[34983] = 8'hd3 ;
            rom[34984] = 8'hfc ;
            rom[34985] = 8'hf5 ;
            rom[34986] = 8'hf6 ;
            rom[34987] = 8'hf8 ;
            rom[34988] = 8'h08 ;
            rom[34989] = 8'h11 ;
            rom[34990] = 8'he5 ;
            rom[34991] = 8'h0f ;
            rom[34992] = 8'h04 ;
            rom[34993] = 8'hd3 ;
            rom[34994] = 8'h0b ;
            rom[34995] = 8'h0f ;
            rom[34996] = 8'hd8 ;
            rom[34997] = 8'h09 ;
            rom[34998] = 8'hea ;
            rom[34999] = 8'hff ;
            rom[35000] = 8'h05 ;
            rom[35001] = 8'hfc ;
            rom[35002] = 8'h0b ;
            rom[35003] = 8'hfe ;
            rom[35004] = 8'h26 ;
            rom[35005] = 8'h13 ;
            rom[35006] = 8'h02 ;
            rom[35007] = 8'hf4 ;
            rom[35008] = 8'hdc ;
            rom[35009] = 8'hfb ;
            rom[35010] = 8'hf3 ;
            rom[35011] = 8'hc4 ;
            rom[35012] = 8'h10 ;
            rom[35013] = 8'h23 ;
            rom[35014] = 8'hef ;
            rom[35015] = 8'h0e ;
            rom[35016] = 8'hef ;
            rom[35017] = 8'h12 ;
            rom[35018] = 8'h0b ;
            rom[35019] = 8'hf5 ;
            rom[35020] = 8'hca ;
            rom[35021] = 8'hfa ;
            rom[35022] = 8'hec ;
            rom[35023] = 8'hdf ;
            rom[35024] = 8'he9 ;
            rom[35025] = 8'hfe ;
            rom[35026] = 8'h2a ;
            rom[35027] = 8'hed ;
            rom[35028] = 8'h1a ;
            rom[35029] = 8'hd9 ;
            rom[35030] = 8'hfa ;
            rom[35031] = 8'h16 ;
            rom[35032] = 8'hfb ;
            rom[35033] = 8'hfb ;
            rom[35034] = 8'h1c ;
            rom[35035] = 8'hdf ;
            rom[35036] = 8'h01 ;
            rom[35037] = 8'hd6 ;
            rom[35038] = 8'h09 ;
            rom[35039] = 8'hd4 ;
            rom[35040] = 8'he0 ;
            rom[35041] = 8'h1d ;
            rom[35042] = 8'h0d ;
            rom[35043] = 8'h1e ;
            rom[35044] = 8'he2 ;
            rom[35045] = 8'hc2 ;
            rom[35046] = 8'h20 ;
            rom[35047] = 8'hef ;
            rom[35048] = 8'h1f ;
            rom[35049] = 8'h0b ;
            rom[35050] = 8'hde ;
            rom[35051] = 8'hce ;
            rom[35052] = 8'hd0 ;
            rom[35053] = 8'h0b ;
            rom[35054] = 8'h20 ;
            rom[35055] = 8'hb6 ;
            rom[35056] = 8'h12 ;
            rom[35057] = 8'h1b ;
            rom[35058] = 8'hfa ;
            rom[35059] = 8'h07 ;
            rom[35060] = 8'hdc ;
            rom[35061] = 8'h0d ;
            rom[35062] = 8'h10 ;
            rom[35063] = 8'h1a ;
            rom[35064] = 8'h0a ;
            rom[35065] = 8'hf9 ;
            rom[35066] = 8'hfe ;
            rom[35067] = 8'h06 ;
            rom[35068] = 8'hc0 ;
            rom[35069] = 8'hfe ;
            rom[35070] = 8'h09 ;
            rom[35071] = 8'hf1 ;
            rom[35072] = 8'h07 ;
            rom[35073] = 8'h19 ;
            rom[35074] = 8'h04 ;
            rom[35075] = 8'he5 ;
            rom[35076] = 8'h04 ;
            rom[35077] = 8'h0f ;
            rom[35078] = 8'hef ;
            rom[35079] = 8'h1f ;
            rom[35080] = 8'h10 ;
            rom[35081] = 8'heb ;
            rom[35082] = 8'h18 ;
            rom[35083] = 8'hf1 ;
            rom[35084] = 8'hf7 ;
            rom[35085] = 8'h02 ;
            rom[35086] = 8'h04 ;
            rom[35087] = 8'h0e ;
            rom[35088] = 8'h0c ;
            rom[35089] = 8'hdc ;
            rom[35090] = 8'hed ;
            rom[35091] = 8'h08 ;
            rom[35092] = 8'h0e ;
            rom[35093] = 8'h03 ;
            rom[35094] = 8'he4 ;
            rom[35095] = 8'hee ;
            rom[35096] = 8'hf3 ;
            rom[35097] = 8'hf1 ;
            rom[35098] = 8'h05 ;
            rom[35099] = 8'h0f ;
            rom[35100] = 8'h0b ;
            rom[35101] = 8'he7 ;
            rom[35102] = 8'h04 ;
            rom[35103] = 8'h98 ;
            rom[35104] = 8'hfa ;
            rom[35105] = 8'hf9 ;
            rom[35106] = 8'hf4 ;
            rom[35107] = 8'h10 ;
            rom[35108] = 8'h08 ;
            rom[35109] = 8'h0f ;
            rom[35110] = 8'hee ;
            rom[35111] = 8'hef ;
            rom[35112] = 8'h0f ;
            rom[35113] = 8'he3 ;
            rom[35114] = 8'h1d ;
            rom[35115] = 8'hf7 ;
            rom[35116] = 8'hf0 ;
            rom[35117] = 8'h18 ;
            rom[35118] = 8'hfe ;
            rom[35119] = 8'hf3 ;
            rom[35120] = 8'hc1 ;
            rom[35121] = 8'hce ;
            rom[35122] = 8'h07 ;
            rom[35123] = 8'hdc ;
            rom[35124] = 8'he2 ;
            rom[35125] = 8'h05 ;
            rom[35126] = 8'hf4 ;
            rom[35127] = 8'hff ;
            rom[35128] = 8'h05 ;
            rom[35129] = 8'he9 ;
            rom[35130] = 8'hfd ;
            rom[35131] = 8'h24 ;
            rom[35132] = 8'he4 ;
            rom[35133] = 8'h15 ;
            rom[35134] = 8'hd7 ;
            rom[35135] = 8'he9 ;
            rom[35136] = 8'h07 ;
            rom[35137] = 8'h17 ;
            rom[35138] = 8'hd3 ;
            rom[35139] = 8'hf2 ;
            rom[35140] = 8'hf1 ;
            rom[35141] = 8'hff ;
            rom[35142] = 8'hea ;
            rom[35143] = 8'hd9 ;
            rom[35144] = 8'h09 ;
            rom[35145] = 8'hfd ;
            rom[35146] = 8'he3 ;
            rom[35147] = 8'hf7 ;
            rom[35148] = 8'hfd ;
            rom[35149] = 8'h0e ;
            rom[35150] = 8'h16 ;
            rom[35151] = 8'h02 ;
            rom[35152] = 8'hfd ;
            rom[35153] = 8'hef ;
            rom[35154] = 8'h1c ;
            rom[35155] = 8'hf0 ;
            rom[35156] = 8'h31 ;
            rom[35157] = 8'hbb ;
            rom[35158] = 8'h1d ;
            rom[35159] = 8'he0 ;
            rom[35160] = 8'hea ;
            rom[35161] = 8'h11 ;
            rom[35162] = 8'hfa ;
            rom[35163] = 8'hf3 ;
            rom[35164] = 8'hcb ;
            rom[35165] = 8'h07 ;
            rom[35166] = 8'he9 ;
            rom[35167] = 8'h04 ;
            rom[35168] = 8'h0a ;
            rom[35169] = 8'h2b ;
            rom[35170] = 8'hf0 ;
            rom[35171] = 8'h0e ;
            rom[35172] = 8'h07 ;
            rom[35173] = 8'hed ;
            rom[35174] = 8'hfc ;
            rom[35175] = 8'hec ;
            rom[35176] = 8'h0d ;
            rom[35177] = 8'heb ;
            rom[35178] = 8'he8 ;
            rom[35179] = 8'hf9 ;
            rom[35180] = 8'h07 ;
            rom[35181] = 8'h1b ;
            rom[35182] = 8'hff ;
            rom[35183] = 8'he9 ;
            rom[35184] = 8'he4 ;
            rom[35185] = 8'hfa ;
            rom[35186] = 8'h13 ;
            rom[35187] = 8'h21 ;
            rom[35188] = 8'hf7 ;
            rom[35189] = 8'h24 ;
            rom[35190] = 8'hec ;
            rom[35191] = 8'hff ;
            rom[35192] = 8'h1a ;
            rom[35193] = 8'h03 ;
            rom[35194] = 8'hf7 ;
            rom[35195] = 8'hdb ;
            rom[35196] = 8'he9 ;
            rom[35197] = 8'h0c ;
            rom[35198] = 8'h14 ;
            rom[35199] = 8'h0c ;
            rom[35200] = 8'hfe ;
            rom[35201] = 8'h0e ;
            rom[35202] = 8'heb ;
            rom[35203] = 8'h1c ;
            rom[35204] = 8'hc8 ;
            rom[35205] = 8'h04 ;
            rom[35206] = 8'h03 ;
            rom[35207] = 8'h19 ;
            rom[35208] = 8'hec ;
            rom[35209] = 8'h18 ;
            rom[35210] = 8'hd8 ;
            rom[35211] = 8'hf9 ;
            rom[35212] = 8'h0e ;
            rom[35213] = 8'he7 ;
            rom[35214] = 8'he2 ;
            rom[35215] = 8'h1f ;
            rom[35216] = 8'hd5 ;
            rom[35217] = 8'hfd ;
            rom[35218] = 8'hf6 ;
            rom[35219] = 8'heb ;
            rom[35220] = 8'h07 ;
            rom[35221] = 8'h02 ;
            rom[35222] = 8'hff ;
            rom[35223] = 8'h0c ;
            rom[35224] = 8'h10 ;
            rom[35225] = 8'hf8 ;
            rom[35226] = 8'hf4 ;
            rom[35227] = 8'h07 ;
            rom[35228] = 8'hf2 ;
            rom[35229] = 8'hdd ;
            rom[35230] = 8'h0b ;
            rom[35231] = 8'h23 ;
            rom[35232] = 8'hf0 ;
            rom[35233] = 8'hd4 ;
            rom[35234] = 8'he5 ;
            rom[35235] = 8'h11 ;
            rom[35236] = 8'h0e ;
            rom[35237] = 8'h0a ;
            rom[35238] = 8'hf5 ;
            rom[35239] = 8'h09 ;
            rom[35240] = 8'hfd ;
            rom[35241] = 8'h10 ;
            rom[35242] = 8'h30 ;
            rom[35243] = 8'h26 ;
            rom[35244] = 8'hfe ;
            rom[35245] = 8'hed ;
            rom[35246] = 8'hd9 ;
            rom[35247] = 8'hfc ;
            rom[35248] = 8'h0e ;
            rom[35249] = 8'hed ;
            rom[35250] = 8'hd1 ;
            rom[35251] = 8'h15 ;
            rom[35252] = 8'h04 ;
            rom[35253] = 8'hf6 ;
            rom[35254] = 8'h0e ;
            rom[35255] = 8'h09 ;
            rom[35256] = 8'he7 ;
            rom[35257] = 8'h02 ;
            rom[35258] = 8'hde ;
            rom[35259] = 8'h00 ;
            rom[35260] = 8'hf1 ;
            rom[35261] = 8'h1a ;
            rom[35262] = 8'h1b ;
            rom[35263] = 8'h0d ;
            rom[35264] = 8'he6 ;
            rom[35265] = 8'hf8 ;
            rom[35266] = 8'h03 ;
            rom[35267] = 8'he7 ;
            rom[35268] = 8'h0f ;
            rom[35269] = 8'h1f ;
            rom[35270] = 8'h0e ;
            rom[35271] = 8'h0d ;
            rom[35272] = 8'hfe ;
            rom[35273] = 8'h01 ;
            rom[35274] = 8'hfd ;
            rom[35275] = 8'hfd ;
            rom[35276] = 8'h09 ;
            rom[35277] = 8'hf9 ;
            rom[35278] = 8'h02 ;
            rom[35279] = 8'h1c ;
            rom[35280] = 8'h22 ;
            rom[35281] = 8'h13 ;
            rom[35282] = 8'h0c ;
            rom[35283] = 8'h02 ;
            rom[35284] = 8'hd1 ;
            rom[35285] = 8'he6 ;
            rom[35286] = 8'h1b ;
            rom[35287] = 8'hef ;
            rom[35288] = 8'hf8 ;
            rom[35289] = 8'h0b ;
            rom[35290] = 8'h14 ;
            rom[35291] = 8'h05 ;
            rom[35292] = 8'h12 ;
            rom[35293] = 8'he1 ;
            rom[35294] = 8'h1a ;
            rom[35295] = 8'hd1 ;
            rom[35296] = 8'heb ;
            rom[35297] = 8'hf8 ;
            rom[35298] = 8'hf5 ;
            rom[35299] = 8'hee ;
            rom[35300] = 8'hfc ;
            rom[35301] = 8'hf2 ;
            rom[35302] = 8'h1b ;
            rom[35303] = 8'h0d ;
            rom[35304] = 8'h02 ;
            rom[35305] = 8'h14 ;
            rom[35306] = 8'h0a ;
            rom[35307] = 8'h03 ;
            rom[35308] = 8'h0d ;
            rom[35309] = 8'he2 ;
            rom[35310] = 8'hde ;
            rom[35311] = 8'h10 ;
            rom[35312] = 8'h06 ;
            rom[35313] = 8'hff ;
            rom[35314] = 8'h05 ;
            rom[35315] = 8'h0b ;
            rom[35316] = 8'h1c ;
            rom[35317] = 8'h0c ;
            rom[35318] = 8'h05 ;
            rom[35319] = 8'hfc ;
            rom[35320] = 8'h0d ;
            rom[35321] = 8'h03 ;
            rom[35322] = 8'h1d ;
            rom[35323] = 8'h19 ;
            rom[35324] = 8'h15 ;
            rom[35325] = 8'h07 ;
            rom[35326] = 8'hfd ;
            rom[35327] = 8'hea ;
            rom[35328] = 8'h18 ;
            rom[35329] = 8'h04 ;
            rom[35330] = 8'hfa ;
            rom[35331] = 8'h14 ;
            rom[35332] = 8'h11 ;
            rom[35333] = 8'hef ;
            rom[35334] = 8'hef ;
            rom[35335] = 8'h0c ;
            rom[35336] = 8'h19 ;
            rom[35337] = 8'h1a ;
            rom[35338] = 8'h01 ;
            rom[35339] = 8'hee ;
            rom[35340] = 8'hd8 ;
            rom[35341] = 8'hcf ;
            rom[35342] = 8'h06 ;
            rom[35343] = 8'he9 ;
            rom[35344] = 8'h1e ;
            rom[35345] = 8'h00 ;
            rom[35346] = 8'h01 ;
            rom[35347] = 8'hfa ;
            rom[35348] = 8'hef ;
            rom[35349] = 8'hee ;
            rom[35350] = 8'hde ;
            rom[35351] = 8'h0a ;
            rom[35352] = 8'hde ;
            rom[35353] = 8'hef ;
            rom[35354] = 8'h0c ;
            rom[35355] = 8'hd7 ;
            rom[35356] = 8'hf6 ;
            rom[35357] = 8'heb ;
            rom[35358] = 8'h11 ;
            rom[35359] = 8'h17 ;
            rom[35360] = 8'hd8 ;
            rom[35361] = 8'h19 ;
            rom[35362] = 8'he7 ;
            rom[35363] = 8'hfa ;
            rom[35364] = 8'hf6 ;
            rom[35365] = 8'hf8 ;
            rom[35366] = 8'hd8 ;
            rom[35367] = 8'hfd ;
            rom[35368] = 8'hf5 ;
            rom[35369] = 8'h16 ;
            rom[35370] = 8'hf9 ;
            rom[35371] = 8'hde ;
            rom[35372] = 8'h1d ;
            rom[35373] = 8'h0d ;
            rom[35374] = 8'h19 ;
            rom[35375] = 8'h0f ;
            rom[35376] = 8'h0c ;
            rom[35377] = 8'h05 ;
            rom[35378] = 8'hf3 ;
            rom[35379] = 8'hfc ;
            rom[35380] = 8'h20 ;
            rom[35381] = 8'hf5 ;
            rom[35382] = 8'he7 ;
            rom[35383] = 8'hf1 ;
            rom[35384] = 8'hf7 ;
            rom[35385] = 8'hf7 ;
            rom[35386] = 8'h0a ;
            rom[35387] = 8'h06 ;
            rom[35388] = 8'h02 ;
            rom[35389] = 8'hf7 ;
            rom[35390] = 8'he3 ;
            rom[35391] = 8'he3 ;
            rom[35392] = 8'hf0 ;
            rom[35393] = 8'he4 ;
            rom[35394] = 8'h03 ;
            rom[35395] = 8'hfc ;
            rom[35396] = 8'h07 ;
            rom[35397] = 8'hfe ;
            rom[35398] = 8'hf7 ;
            rom[35399] = 8'hff ;
            rom[35400] = 8'hfa ;
            rom[35401] = 8'hd2 ;
            rom[35402] = 8'h08 ;
            rom[35403] = 8'hfb ;
            rom[35404] = 8'h0c ;
            rom[35405] = 8'hf7 ;
            rom[35406] = 8'hcf ;
            rom[35407] = 8'hf9 ;
            rom[35408] = 8'hf8 ;
            rom[35409] = 8'hbc ;
            rom[35410] = 8'hed ;
            rom[35411] = 8'h00 ;
            rom[35412] = 8'hfe ;
            rom[35413] = 8'h0a ;
            rom[35414] = 8'hda ;
            rom[35415] = 8'hff ;
            rom[35416] = 8'h1a ;
            rom[35417] = 8'hf2 ;
            rom[35418] = 8'h1a ;
            rom[35419] = 8'h13 ;
            rom[35420] = 8'h07 ;
            rom[35421] = 8'h05 ;
            rom[35422] = 8'h03 ;
            rom[35423] = 8'h18 ;
            rom[35424] = 8'hf1 ;
            rom[35425] = 8'hc1 ;
            rom[35426] = 8'hfb ;
            rom[35427] = 8'hcc ;
            rom[35428] = 8'hd8 ;
            rom[35429] = 8'he9 ;
            rom[35430] = 8'hfa ;
            rom[35431] = 8'hfc ;
            rom[35432] = 8'hb1 ;
            rom[35433] = 8'h9f ;
            rom[35434] = 8'he7 ;
            rom[35435] = 8'h21 ;
            rom[35436] = 8'h0a ;
            rom[35437] = 8'hee ;
            rom[35438] = 8'h05 ;
            rom[35439] = 8'hfc ;
            rom[35440] = 8'hef ;
            rom[35441] = 8'h10 ;
            rom[35442] = 8'h1b ;
            rom[35443] = 8'hdb ;
            rom[35444] = 8'hf8 ;
            rom[35445] = 8'h0a ;
            rom[35446] = 8'hfd ;
            rom[35447] = 8'he9 ;
            rom[35448] = 8'hf6 ;
            rom[35449] = 8'hdf ;
            rom[35450] = 8'h13 ;
            rom[35451] = 8'h09 ;
            rom[35452] = 8'h14 ;
            rom[35453] = 8'he3 ;
            rom[35454] = 8'hf8 ;
            rom[35455] = 8'hed ;
            rom[35456] = 8'he4 ;
            rom[35457] = 8'hf3 ;
            rom[35458] = 8'h19 ;
            rom[35459] = 8'h02 ;
            rom[35460] = 8'hff ;
            rom[35461] = 8'hfe ;
            rom[35462] = 8'h15 ;
            rom[35463] = 8'he0 ;
            rom[35464] = 8'hf7 ;
            rom[35465] = 8'hee ;
            rom[35466] = 8'h17 ;
            rom[35467] = 8'h0e ;
            rom[35468] = 8'h09 ;
            rom[35469] = 8'hfe ;
            rom[35470] = 8'h07 ;
            rom[35471] = 8'hf1 ;
            rom[35472] = 8'hc6 ;
            rom[35473] = 8'heb ;
            rom[35474] = 8'h13 ;
            rom[35475] = 8'hde ;
            rom[35476] = 8'h0b ;
            rom[35477] = 8'h16 ;
            rom[35478] = 8'h02 ;
            rom[35479] = 8'hff ;
            rom[35480] = 8'h16 ;
            rom[35481] = 8'hf7 ;
            rom[35482] = 8'h04 ;
            rom[35483] = 8'he9 ;
            rom[35484] = 8'hfd ;
            rom[35485] = 8'h18 ;
            rom[35486] = 8'hf7 ;
            rom[35487] = 8'h0a ;
            rom[35488] = 8'he5 ;
            rom[35489] = 8'ha8 ;
            rom[35490] = 8'he6 ;
            rom[35491] = 8'h1c ;
            rom[35492] = 8'hfc ;
            rom[35493] = 8'hf0 ;
            rom[35494] = 8'h26 ;
            rom[35495] = 8'h16 ;
            rom[35496] = 8'h07 ;
            rom[35497] = 8'hf0 ;
            rom[35498] = 8'he4 ;
            rom[35499] = 8'h03 ;
            rom[35500] = 8'h14 ;
            rom[35501] = 8'hfa ;
            rom[35502] = 8'h0f ;
            rom[35503] = 8'hd4 ;
            rom[35504] = 8'hf3 ;
            rom[35505] = 8'hef ;
            rom[35506] = 8'h23 ;
            rom[35507] = 8'hcc ;
            rom[35508] = 8'h09 ;
            rom[35509] = 8'h07 ;
            rom[35510] = 8'h0a ;
            rom[35511] = 8'hd3 ;
            rom[35512] = 8'hf6 ;
            rom[35513] = 8'hf7 ;
            rom[35514] = 8'h18 ;
            rom[35515] = 8'h25 ;
            rom[35516] = 8'he8 ;
            rom[35517] = 8'hc6 ;
            rom[35518] = 8'hf1 ;
            rom[35519] = 8'hcd ;
            rom[35520] = 8'h28 ;
            rom[35521] = 8'h0f ;
            rom[35522] = 8'hf4 ;
            rom[35523] = 8'he3 ;
            rom[35524] = 8'h22 ;
            rom[35525] = 8'h0f ;
            rom[35526] = 8'hba ;
            rom[35527] = 8'h1a ;
            rom[35528] = 8'hd1 ;
            rom[35529] = 8'h03 ;
            rom[35530] = 8'h08 ;
            rom[35531] = 8'h07 ;
            rom[35532] = 8'hf2 ;
            rom[35533] = 8'he0 ;
            rom[35534] = 8'hcf ;
            rom[35535] = 8'hec ;
            rom[35536] = 8'hfe ;
            rom[35537] = 8'hfb ;
            rom[35538] = 8'h0b ;
            rom[35539] = 8'h0c ;
            rom[35540] = 8'hb7 ;
            rom[35541] = 8'hfe ;
            rom[35542] = 8'he3 ;
            rom[35543] = 8'he4 ;
            rom[35544] = 8'h01 ;
            rom[35545] = 8'hf2 ;
            rom[35546] = 8'he8 ;
            rom[35547] = 8'hf9 ;
            rom[35548] = 8'h13 ;
            rom[35549] = 8'hea ;
            rom[35550] = 8'hff ;
            rom[35551] = 8'hf8 ;
            rom[35552] = 8'hd6 ;
            rom[35553] = 8'he2 ;
            rom[35554] = 8'hf3 ;
            rom[35555] = 8'hf9 ;
            rom[35556] = 8'h19 ;
            rom[35557] = 8'h09 ;
            rom[35558] = 8'hfe ;
            rom[35559] = 8'hbf ;
            rom[35560] = 8'h20 ;
            rom[35561] = 8'hf0 ;
            rom[35562] = 8'hf3 ;
            rom[35563] = 8'h2a ;
            rom[35564] = 8'hc5 ;
            rom[35565] = 8'h32 ;
            rom[35566] = 8'hf1 ;
            rom[35567] = 8'h12 ;
            rom[35568] = 8'h01 ;
            rom[35569] = 8'hf0 ;
            rom[35570] = 8'h04 ;
            rom[35571] = 8'hf1 ;
            rom[35572] = 8'h05 ;
            rom[35573] = 8'hfc ;
            rom[35574] = 8'h04 ;
            rom[35575] = 8'heb ;
            rom[35576] = 8'hf0 ;
            rom[35577] = 8'h18 ;
            rom[35578] = 8'h0e ;
            rom[35579] = 8'hf8 ;
            rom[35580] = 8'h00 ;
            rom[35581] = 8'h10 ;
            rom[35582] = 8'hef ;
            rom[35583] = 8'hfa ;
            rom[35584] = 8'h23 ;
            rom[35585] = 8'hf9 ;
            rom[35586] = 8'h15 ;
            rom[35587] = 8'hf3 ;
            rom[35588] = 8'h0a ;
            rom[35589] = 8'hf8 ;
            rom[35590] = 8'hf1 ;
            rom[35591] = 8'hff ;
            rom[35592] = 8'hff ;
            rom[35593] = 8'hf9 ;
            rom[35594] = 8'he6 ;
            rom[35595] = 8'hfd ;
            rom[35596] = 8'hcd ;
            rom[35597] = 8'h13 ;
            rom[35598] = 8'hcc ;
            rom[35599] = 8'h00 ;
            rom[35600] = 8'h1e ;
            rom[35601] = 8'h07 ;
            rom[35602] = 8'h01 ;
            rom[35603] = 8'h15 ;
            rom[35604] = 8'hf7 ;
            rom[35605] = 8'h00 ;
            rom[35606] = 8'hfa ;
            rom[35607] = 8'hdd ;
            rom[35608] = 8'hff ;
            rom[35609] = 8'h0f ;
            rom[35610] = 8'hff ;
            rom[35611] = 8'h08 ;
            rom[35612] = 8'h06 ;
            rom[35613] = 8'h28 ;
            rom[35614] = 8'h0f ;
            rom[35615] = 8'hf4 ;
            rom[35616] = 8'he1 ;
            rom[35617] = 8'h20 ;
            rom[35618] = 8'hff ;
            rom[35619] = 8'hf1 ;
            rom[35620] = 8'h0a ;
            rom[35621] = 8'he8 ;
            rom[35622] = 8'h0a ;
            rom[35623] = 8'h05 ;
            rom[35624] = 8'hd6 ;
            rom[35625] = 8'hf5 ;
            rom[35626] = 8'h0a ;
            rom[35627] = 8'he6 ;
            rom[35628] = 8'hed ;
            rom[35629] = 8'hf5 ;
            rom[35630] = 8'he8 ;
            rom[35631] = 8'he6 ;
            rom[35632] = 8'he5 ;
            rom[35633] = 8'h19 ;
            rom[35634] = 8'h09 ;
            rom[35635] = 8'hfb ;
            rom[35636] = 8'hdd ;
            rom[35637] = 8'hd8 ;
            rom[35638] = 8'hfd ;
            rom[35639] = 8'h08 ;
            rom[35640] = 8'hfa ;
            rom[35641] = 8'h09 ;
            rom[35642] = 8'h05 ;
            rom[35643] = 8'he7 ;
            rom[35644] = 8'hef ;
            rom[35645] = 8'h0c ;
            rom[35646] = 8'hf1 ;
            rom[35647] = 8'he5 ;
            rom[35648] = 8'hff ;
            rom[35649] = 8'hf8 ;
            rom[35650] = 8'hfc ;
            rom[35651] = 8'hfa ;
            rom[35652] = 8'h15 ;
            rom[35653] = 8'hf8 ;
            rom[35654] = 8'h07 ;
            rom[35655] = 8'h02 ;
            rom[35656] = 8'h1c ;
            rom[35657] = 8'hf7 ;
            rom[35658] = 8'hf2 ;
            rom[35659] = 8'hea ;
            rom[35660] = 8'h01 ;
            rom[35661] = 8'h0e ;
            rom[35662] = 8'he8 ;
            rom[35663] = 8'hdd ;
            rom[35664] = 8'hf2 ;
            rom[35665] = 8'hd5 ;
            rom[35666] = 8'hf2 ;
            rom[35667] = 8'h06 ;
            rom[35668] = 8'h08 ;
            rom[35669] = 8'heb ;
            rom[35670] = 8'h0e ;
            rom[35671] = 8'h13 ;
            rom[35672] = 8'he1 ;
            rom[35673] = 8'he8 ;
            rom[35674] = 8'hd8 ;
            rom[35675] = 8'hb4 ;
            rom[35676] = 8'hf3 ;
            rom[35677] = 8'h0f ;
            rom[35678] = 8'hf2 ;
            rom[35679] = 8'hdc ;
            rom[35680] = 8'h04 ;
            rom[35681] = 8'hd7 ;
            rom[35682] = 8'hc3 ;
            rom[35683] = 8'h29 ;
            rom[35684] = 8'h0c ;
            rom[35685] = 8'hf9 ;
            rom[35686] = 8'hff ;
            rom[35687] = 8'h09 ;
            rom[35688] = 8'hd5 ;
            rom[35689] = 8'heb ;
            rom[35690] = 8'hf8 ;
            rom[35691] = 8'h01 ;
            rom[35692] = 8'he1 ;
            rom[35693] = 8'hf6 ;
            rom[35694] = 8'hed ;
            rom[35695] = 8'hf0 ;
            rom[35696] = 8'hfc ;
            rom[35697] = 8'he0 ;
            rom[35698] = 8'h17 ;
            rom[35699] = 8'hfa ;
            rom[35700] = 8'hd0 ;
            rom[35701] = 8'hfb ;
            rom[35702] = 8'hc9 ;
            rom[35703] = 8'hd6 ;
            rom[35704] = 8'hff ;
            rom[35705] = 8'hf5 ;
            rom[35706] = 8'hcf ;
            rom[35707] = 8'hf0 ;
            rom[35708] = 8'he8 ;
            rom[35709] = 8'hf8 ;
            rom[35710] = 8'h08 ;
            rom[35711] = 8'hfa ;
            rom[35712] = 8'h0f ;
            rom[35713] = 8'h00 ;
            rom[35714] = 8'hf0 ;
            rom[35715] = 8'h01 ;
            rom[35716] = 8'h03 ;
            rom[35717] = 8'hdf ;
            rom[35718] = 8'h19 ;
            rom[35719] = 8'hff ;
            rom[35720] = 8'hfd ;
            rom[35721] = 8'h09 ;
            rom[35722] = 8'hcd ;
            rom[35723] = 8'hee ;
            rom[35724] = 8'hfc ;
            rom[35725] = 8'h31 ;
            rom[35726] = 8'hd5 ;
            rom[35727] = 8'hfb ;
            rom[35728] = 8'h05 ;
            rom[35729] = 8'he7 ;
            rom[35730] = 8'h18 ;
            rom[35731] = 8'h00 ;
            rom[35732] = 8'h16 ;
            rom[35733] = 8'hc9 ;
            rom[35734] = 8'h25 ;
            rom[35735] = 8'hfa ;
            rom[35736] = 8'hf2 ;
            rom[35737] = 8'h19 ;
            rom[35738] = 8'hd8 ;
            rom[35739] = 8'h02 ;
            rom[35740] = 8'h0a ;
            rom[35741] = 8'h1d ;
            rom[35742] = 8'hf8 ;
            rom[35743] = 8'hf4 ;
            rom[35744] = 8'hee ;
            rom[35745] = 8'he2 ;
            rom[35746] = 8'hf5 ;
            rom[35747] = 8'h12 ;
            rom[35748] = 8'hfa ;
            rom[35749] = 8'hd4 ;
            rom[35750] = 8'h0f ;
            rom[35751] = 8'hd4 ;
            rom[35752] = 8'hf0 ;
            rom[35753] = 8'hde ;
            rom[35754] = 8'h19 ;
            rom[35755] = 8'hc7 ;
            rom[35756] = 8'h00 ;
            rom[35757] = 8'hf4 ;
            rom[35758] = 8'hde ;
            rom[35759] = 8'h21 ;
            rom[35760] = 8'hfe ;
            rom[35761] = 8'h0e ;
            rom[35762] = 8'h19 ;
            rom[35763] = 8'h16 ;
            rom[35764] = 8'hf6 ;
            rom[35765] = 8'hf6 ;
            rom[35766] = 8'h01 ;
            rom[35767] = 8'hf0 ;
            rom[35768] = 8'heb ;
            rom[35769] = 8'h0c ;
            rom[35770] = 8'hec ;
            rom[35771] = 8'hf8 ;
            rom[35772] = 8'hf6 ;
            rom[35773] = 8'hfb ;
            rom[35774] = 8'he9 ;
            rom[35775] = 8'h13 ;
            rom[35776] = 8'he9 ;
            rom[35777] = 8'hfe ;
            rom[35778] = 8'h05 ;
            rom[35779] = 8'hfd ;
            rom[35780] = 8'he9 ;
            rom[35781] = 8'h18 ;
            rom[35782] = 8'hfd ;
            rom[35783] = 8'h0f ;
            rom[35784] = 8'hf4 ;
            rom[35785] = 8'h0c ;
            rom[35786] = 8'h0e ;
            rom[35787] = 8'h03 ;
            rom[35788] = 8'hff ;
            rom[35789] = 8'hee ;
            rom[35790] = 8'h0a ;
            rom[35791] = 8'h15 ;
            rom[35792] = 8'h14 ;
            rom[35793] = 8'h0e ;
            rom[35794] = 8'he6 ;
            rom[35795] = 8'h04 ;
            rom[35796] = 8'he0 ;
            rom[35797] = 8'h0a ;
            rom[35798] = 8'hec ;
            rom[35799] = 8'h07 ;
            rom[35800] = 8'hfb ;
            rom[35801] = 8'hdf ;
            rom[35802] = 8'hfe ;
            rom[35803] = 8'hf5 ;
            rom[35804] = 8'hd9 ;
            rom[35805] = 8'hf3 ;
            rom[35806] = 8'h05 ;
            rom[35807] = 8'hf6 ;
            rom[35808] = 8'h05 ;
            rom[35809] = 8'h2f ;
            rom[35810] = 8'hee ;
            rom[35811] = 8'h19 ;
            rom[35812] = 8'hfe ;
            rom[35813] = 8'h1b ;
            rom[35814] = 8'h0a ;
            rom[35815] = 8'h0f ;
            rom[35816] = 8'hfb ;
            rom[35817] = 8'h0f ;
            rom[35818] = 8'hf1 ;
            rom[35819] = 8'h20 ;
            rom[35820] = 8'he0 ;
            rom[35821] = 8'h0e ;
            rom[35822] = 8'hc8 ;
            rom[35823] = 8'hc4 ;
            rom[35824] = 8'hfd ;
            rom[35825] = 8'he7 ;
            rom[35826] = 8'h01 ;
            rom[35827] = 8'hd6 ;
            rom[35828] = 8'h17 ;
            rom[35829] = 8'hfa ;
            rom[35830] = 8'hf9 ;
            rom[35831] = 8'hf0 ;
            rom[35832] = 8'h2d ;
            rom[35833] = 8'hf0 ;
            rom[35834] = 8'hfe ;
            rom[35835] = 8'h1e ;
            rom[35836] = 8'hea ;
            rom[35837] = 8'hf6 ;
            rom[35838] = 8'hf3 ;
            rom[35839] = 8'h05 ;
            rom[35840] = 8'hd0 ;
            rom[35841] = 8'h12 ;
            rom[35842] = 8'hf2 ;
            rom[35843] = 8'hda ;
            rom[35844] = 8'hfa ;
            rom[35845] = 8'he5 ;
            rom[35846] = 8'h0a ;
            rom[35847] = 8'hfb ;
            rom[35848] = 8'h00 ;
            rom[35849] = 8'hed ;
            rom[35850] = 8'h09 ;
            rom[35851] = 8'h0c ;
            rom[35852] = 8'h06 ;
            rom[35853] = 8'hdb ;
            rom[35854] = 8'hfe ;
            rom[35855] = 8'h29 ;
            rom[35856] = 8'he5 ;
            rom[35857] = 8'hd5 ;
            rom[35858] = 8'hfc ;
            rom[35859] = 8'h17 ;
            rom[35860] = 8'h14 ;
            rom[35861] = 8'h17 ;
            rom[35862] = 8'hee ;
            rom[35863] = 8'h11 ;
            rom[35864] = 8'h16 ;
            rom[35865] = 8'hf4 ;
            rom[35866] = 8'hea ;
            rom[35867] = 8'h05 ;
            rom[35868] = 8'hcc ;
            rom[35869] = 8'h03 ;
            rom[35870] = 8'hf2 ;
            rom[35871] = 8'hdc ;
            rom[35872] = 8'h24 ;
            rom[35873] = 8'hd1 ;
            rom[35874] = 8'he5 ;
            rom[35875] = 8'hf4 ;
            rom[35876] = 8'h16 ;
            rom[35877] = 8'h33 ;
            rom[35878] = 8'h11 ;
            rom[35879] = 8'hfc ;
            rom[35880] = 8'hff ;
            rom[35881] = 8'he2 ;
            rom[35882] = 8'hf0 ;
            rom[35883] = 8'h18 ;
            rom[35884] = 8'h08 ;
            rom[35885] = 8'hfe ;
            rom[35886] = 8'h0e ;
            rom[35887] = 8'hd8 ;
            rom[35888] = 8'hf2 ;
            rom[35889] = 8'hf7 ;
            rom[35890] = 8'hfc ;
            rom[35891] = 8'hfe ;
            rom[35892] = 8'hd7 ;
            rom[35893] = 8'hf3 ;
            rom[35894] = 8'hf5 ;
            rom[35895] = 8'hf6 ;
            rom[35896] = 8'h21 ;
            rom[35897] = 8'hf8 ;
            rom[35898] = 8'h17 ;
            rom[35899] = 8'hf5 ;
            rom[35900] = 8'h1d ;
            rom[35901] = 8'h1d ;
            rom[35902] = 8'h07 ;
            rom[35903] = 8'h02 ;
            rom[35904] = 8'h0c ;
            rom[35905] = 8'h0e ;
            rom[35906] = 8'hff ;
            rom[35907] = 8'hfd ;
            rom[35908] = 8'hd4 ;
            rom[35909] = 8'h08 ;
            rom[35910] = 8'he0 ;
            rom[35911] = 8'hf7 ;
            rom[35912] = 8'hc8 ;
            rom[35913] = 8'hfe ;
            rom[35914] = 8'hfe ;
            rom[35915] = 8'hfb ;
            rom[35916] = 8'hc1 ;
            rom[35917] = 8'hfd ;
            rom[35918] = 8'h0f ;
            rom[35919] = 8'h25 ;
            rom[35920] = 8'h2e ;
            rom[35921] = 8'h0f ;
            rom[35922] = 8'h22 ;
            rom[35923] = 8'hf3 ;
            rom[35924] = 8'h27 ;
            rom[35925] = 8'hde ;
            rom[35926] = 8'hfc ;
            rom[35927] = 8'hca ;
            rom[35928] = 8'hdc ;
            rom[35929] = 8'h0b ;
            rom[35930] = 8'h05 ;
            rom[35931] = 8'he6 ;
            rom[35932] = 8'he2 ;
            rom[35933] = 8'h04 ;
            rom[35934] = 8'h1b ;
            rom[35935] = 8'hf8 ;
            rom[35936] = 8'hfc ;
            rom[35937] = 8'h08 ;
            rom[35938] = 8'hfa ;
            rom[35939] = 8'h23 ;
            rom[35940] = 8'h06 ;
            rom[35941] = 8'hf7 ;
            rom[35942] = 8'h09 ;
            rom[35943] = 8'hec ;
            rom[35944] = 8'h0a ;
            rom[35945] = 8'hfa ;
            rom[35946] = 8'hf9 ;
            rom[35947] = 8'h0e ;
            rom[35948] = 8'he6 ;
            rom[35949] = 8'h0d ;
            rom[35950] = 8'hee ;
            rom[35951] = 8'h0a ;
            rom[35952] = 8'hff ;
            rom[35953] = 8'hf1 ;
            rom[35954] = 8'hf9 ;
            rom[35955] = 8'h28 ;
            rom[35956] = 8'h32 ;
            rom[35957] = 8'h26 ;
            rom[35958] = 8'h13 ;
            rom[35959] = 8'h06 ;
            rom[35960] = 8'h03 ;
            rom[35961] = 8'h12 ;
            rom[35962] = 8'hf3 ;
            rom[35963] = 8'hec ;
            rom[35964] = 8'h08 ;
            rom[35965] = 8'hf6 ;
            rom[35966] = 8'hff ;
            rom[35967] = 8'h0b ;
            rom[35968] = 8'hcc ;
            rom[35969] = 8'h10 ;
            rom[35970] = 8'h09 ;
            rom[35971] = 8'hd7 ;
            rom[35972] = 8'hd5 ;
            rom[35973] = 8'h0f ;
            rom[35974] = 8'hee ;
            rom[35975] = 8'hf3 ;
            rom[35976] = 8'h05 ;
            rom[35977] = 8'h08 ;
            rom[35978] = 8'h0c ;
            rom[35979] = 8'h0a ;
            rom[35980] = 8'hd7 ;
            rom[35981] = 8'hfc ;
            rom[35982] = 8'hdf ;
            rom[35983] = 8'h0c ;
            rom[35984] = 8'hf5 ;
            rom[35985] = 8'h05 ;
            rom[35986] = 8'h00 ;
            rom[35987] = 8'hee ;
            rom[35988] = 8'h17 ;
            rom[35989] = 8'h06 ;
            rom[35990] = 8'hfc ;
            rom[35991] = 8'h0d ;
            rom[35992] = 8'he1 ;
            rom[35993] = 8'h26 ;
            rom[35994] = 8'hcb ;
            rom[35995] = 8'h2e ;
            rom[35996] = 8'hef ;
            rom[35997] = 8'h1e ;
            rom[35998] = 8'hf4 ;
            rom[35999] = 8'hf4 ;
            rom[36000] = 8'h1f ;
            rom[36001] = 8'h0d ;
            rom[36002] = 8'h01 ;
            rom[36003] = 8'hfe ;
            rom[36004] = 8'h1e ;
            rom[36005] = 8'h02 ;
            rom[36006] = 8'hd8 ;
            rom[36007] = 8'hf3 ;
            rom[36008] = 8'hc9 ;
            rom[36009] = 8'hd2 ;
            rom[36010] = 8'hf2 ;
            rom[36011] = 8'h1c ;
            rom[36012] = 8'hf4 ;
            rom[36013] = 8'hcb ;
            rom[36014] = 8'hff ;
            rom[36015] = 8'hfb ;
            rom[36016] = 8'hf0 ;
            rom[36017] = 8'h08 ;
            rom[36018] = 8'h00 ;
            rom[36019] = 8'h11 ;
            rom[36020] = 8'h0b ;
            rom[36021] = 8'h1a ;
            rom[36022] = 8'h06 ;
            rom[36023] = 8'hdf ;
            rom[36024] = 8'hdd ;
            rom[36025] = 8'h1a ;
            rom[36026] = 8'hf4 ;
            rom[36027] = 8'hf8 ;
            rom[36028] = 8'h06 ;
            rom[36029] = 8'hd8 ;
            rom[36030] = 8'h13 ;
            rom[36031] = 8'h13 ;
            rom[36032] = 8'hf2 ;
            rom[36033] = 8'hee ;
            rom[36034] = 8'h10 ;
            rom[36035] = 8'h13 ;
            rom[36036] = 8'hcf ;
            rom[36037] = 8'h12 ;
            rom[36038] = 8'h1a ;
            rom[36039] = 8'h07 ;
            rom[36040] = 8'hdc ;
            rom[36041] = 8'h08 ;
            rom[36042] = 8'he9 ;
            rom[36043] = 8'h05 ;
            rom[36044] = 8'hf9 ;
            rom[36045] = 8'hd1 ;
            rom[36046] = 8'h0a ;
            rom[36047] = 8'he6 ;
            rom[36048] = 8'h0d ;
            rom[36049] = 8'hf2 ;
            rom[36050] = 8'h01 ;
            rom[36051] = 8'he9 ;
            rom[36052] = 8'hd4 ;
            rom[36053] = 8'hdf ;
            rom[36054] = 8'hef ;
            rom[36055] = 8'h2e ;
            rom[36056] = 8'h0c ;
            rom[36057] = 8'hee ;
            rom[36058] = 8'h11 ;
            rom[36059] = 8'hdb ;
            rom[36060] = 8'hfd ;
            rom[36061] = 8'heb ;
            rom[36062] = 8'hf1 ;
            rom[36063] = 8'hf7 ;
            rom[36064] = 8'h09 ;
            rom[36065] = 8'hf3 ;
            rom[36066] = 8'hdd ;
            rom[36067] = 8'h14 ;
            rom[36068] = 8'h07 ;
            rom[36069] = 8'h09 ;
            rom[36070] = 8'h07 ;
            rom[36071] = 8'h11 ;
            rom[36072] = 8'hf4 ;
            rom[36073] = 8'hfd ;
            rom[36074] = 8'hf9 ;
            rom[36075] = 8'he1 ;
            rom[36076] = 8'h0d ;
            rom[36077] = 8'h0a ;
            rom[36078] = 8'h0b ;
            rom[36079] = 8'hf7 ;
            rom[36080] = 8'h0c ;
            rom[36081] = 8'h07 ;
            rom[36082] = 8'hf7 ;
            rom[36083] = 8'h1b ;
            rom[36084] = 8'hfe ;
            rom[36085] = 8'hee ;
            rom[36086] = 8'he9 ;
            rom[36087] = 8'h27 ;
            rom[36088] = 8'h04 ;
            rom[36089] = 8'hfb ;
            rom[36090] = 8'hdc ;
            rom[36091] = 8'hf8 ;
            rom[36092] = 8'h12 ;
            rom[36093] = 8'hf0 ;
            rom[36094] = 8'hf2 ;
            rom[36095] = 8'h03 ;
            rom[36096] = 8'hfc ;
            rom[36097] = 8'hf2 ;
            rom[36098] = 8'h0f ;
            rom[36099] = 8'he2 ;
            rom[36100] = 8'hfd ;
            rom[36101] = 8'hf4 ;
            rom[36102] = 8'h20 ;
            rom[36103] = 8'hf7 ;
            rom[36104] = 8'hf6 ;
            rom[36105] = 8'h04 ;
            rom[36106] = 8'h14 ;
            rom[36107] = 8'h33 ;
            rom[36108] = 8'hd3 ;
            rom[36109] = 8'h17 ;
            rom[36110] = 8'h1c ;
            rom[36111] = 8'hfc ;
            rom[36112] = 8'he3 ;
            rom[36113] = 8'h12 ;
            rom[36114] = 8'h20 ;
            rom[36115] = 8'h1b ;
            rom[36116] = 8'h01 ;
            rom[36117] = 8'he8 ;
            rom[36118] = 8'h21 ;
            rom[36119] = 8'h19 ;
            rom[36120] = 8'hf6 ;
            rom[36121] = 8'hd7 ;
            rom[36122] = 8'hfe ;
            rom[36123] = 8'hd8 ;
            rom[36124] = 8'hfe ;
            rom[36125] = 8'hed ;
            rom[36126] = 8'hc5 ;
            rom[36127] = 8'hf4 ;
            rom[36128] = 8'hfd ;
            rom[36129] = 8'h0b ;
            rom[36130] = 8'h08 ;
            rom[36131] = 8'h04 ;
            rom[36132] = 8'h07 ;
            rom[36133] = 8'he3 ;
            rom[36134] = 8'hf2 ;
            rom[36135] = 8'hd4 ;
            rom[36136] = 8'h05 ;
            rom[36137] = 8'he9 ;
            rom[36138] = 8'hec ;
            rom[36139] = 8'hee ;
            rom[36140] = 8'hee ;
            rom[36141] = 8'hef ;
            rom[36142] = 8'h14 ;
            rom[36143] = 8'hdc ;
            rom[36144] = 8'h11 ;
            rom[36145] = 8'hca ;
            rom[36146] = 8'h03 ;
            rom[36147] = 8'hf3 ;
            rom[36148] = 8'he5 ;
            rom[36149] = 8'hf8 ;
            rom[36150] = 8'h19 ;
            rom[36151] = 8'hec ;
            rom[36152] = 8'h17 ;
            rom[36153] = 8'h08 ;
            rom[36154] = 8'hcc ;
            rom[36155] = 8'h2c ;
            rom[36156] = 8'h17 ;
            rom[36157] = 8'h08 ;
            rom[36158] = 8'h1d ;
            rom[36159] = 8'hfb ;
            rom[36160] = 8'hf3 ;
            rom[36161] = 8'h02 ;
            rom[36162] = 8'h0a ;
            rom[36163] = 8'h1c ;
            rom[36164] = 8'hd9 ;
            rom[36165] = 8'h07 ;
            rom[36166] = 8'hc7 ;
            rom[36167] = 8'h1f ;
            rom[36168] = 8'hf4 ;
            rom[36169] = 8'h2f ;
            rom[36170] = 8'h0f ;
            rom[36171] = 8'h0d ;
            rom[36172] = 8'heb ;
            rom[36173] = 8'h2a ;
            rom[36174] = 8'hec ;
            rom[36175] = 8'h11 ;
            rom[36176] = 8'hfe ;
            rom[36177] = 8'h27 ;
            rom[36178] = 8'h0a ;
            rom[36179] = 8'hf9 ;
            rom[36180] = 8'hfe ;
            rom[36181] = 8'h0a ;
            rom[36182] = 8'he8 ;
            rom[36183] = 8'h11 ;
            rom[36184] = 8'hdf ;
            rom[36185] = 8'hff ;
            rom[36186] = 8'hef ;
            rom[36187] = 8'h05 ;
            rom[36188] = 8'hf6 ;
            rom[36189] = 8'hf4 ;
            rom[36190] = 8'h19 ;
            rom[36191] = 8'h0d ;
            rom[36192] = 8'hfc ;
            rom[36193] = 8'he9 ;
            rom[36194] = 8'h2e ;
            rom[36195] = 8'h0e ;
            rom[36196] = 8'hf7 ;
            rom[36197] = 8'h05 ;
            rom[36198] = 8'h06 ;
            rom[36199] = 8'he8 ;
            rom[36200] = 8'h1a ;
            rom[36201] = 8'hed ;
            rom[36202] = 8'he1 ;
            rom[36203] = 8'h10 ;
            rom[36204] = 8'he2 ;
            rom[36205] = 8'hed ;
            rom[36206] = 8'h21 ;
            rom[36207] = 8'h0d ;
            rom[36208] = 8'h00 ;
            rom[36209] = 8'hf1 ;
            rom[36210] = 8'hef ;
            rom[36211] = 8'hf7 ;
            rom[36212] = 8'h14 ;
            rom[36213] = 8'h03 ;
            rom[36214] = 8'h00 ;
            rom[36215] = 8'h01 ;
            rom[36216] = 8'h05 ;
            rom[36217] = 8'h2d ;
            rom[36218] = 8'h09 ;
            rom[36219] = 8'hfd ;
            rom[36220] = 8'h14 ;
            rom[36221] = 8'h19 ;
            rom[36222] = 8'hf8 ;
            rom[36223] = 8'h03 ;
            rom[36224] = 8'h18 ;
            rom[36225] = 8'h0e ;
            rom[36226] = 8'h32 ;
            rom[36227] = 8'h09 ;
            rom[36228] = 8'he8 ;
            rom[36229] = 8'he8 ;
            rom[36230] = 8'hfc ;
            rom[36231] = 8'h08 ;
            rom[36232] = 8'h05 ;
            rom[36233] = 8'hf9 ;
            rom[36234] = 8'h06 ;
            rom[36235] = 8'hd4 ;
            rom[36236] = 8'hc2 ;
            rom[36237] = 8'hf8 ;
            rom[36238] = 8'hfe ;
            rom[36239] = 8'hec ;
            rom[36240] = 8'he7 ;
            rom[36241] = 8'h31 ;
            rom[36242] = 8'h01 ;
            rom[36243] = 8'h06 ;
            rom[36244] = 8'hea ;
            rom[36245] = 8'hf8 ;
            rom[36246] = 8'hec ;
            rom[36247] = 8'hc8 ;
            rom[36248] = 8'hd6 ;
            rom[36249] = 8'h0a ;
            rom[36250] = 8'he1 ;
            rom[36251] = 8'h03 ;
            rom[36252] = 8'h0c ;
            rom[36253] = 8'h09 ;
            rom[36254] = 8'h04 ;
            rom[36255] = 8'h19 ;
            rom[36256] = 8'hed ;
            rom[36257] = 8'h07 ;
            rom[36258] = 8'hf7 ;
            rom[36259] = 8'hf2 ;
            rom[36260] = 8'h0c ;
            rom[36261] = 8'h06 ;
            rom[36262] = 8'hf4 ;
            rom[36263] = 8'h02 ;
            rom[36264] = 8'hcd ;
            rom[36265] = 8'hff ;
            rom[36266] = 8'hef ;
            rom[36267] = 8'h08 ;
            rom[36268] = 8'hda ;
            rom[36269] = 8'hda ;
            rom[36270] = 8'he0 ;
            rom[36271] = 8'hf5 ;
            rom[36272] = 8'h05 ;
            rom[36273] = 8'hf0 ;
            rom[36274] = 8'hd1 ;
            rom[36275] = 8'he6 ;
            rom[36276] = 8'heb ;
            rom[36277] = 8'h07 ;
            rom[36278] = 8'hfc ;
            rom[36279] = 8'hf9 ;
            rom[36280] = 8'hf3 ;
            rom[36281] = 8'h01 ;
            rom[36282] = 8'hf7 ;
            rom[36283] = 8'h1a ;
            rom[36284] = 8'h20 ;
            rom[36285] = 8'he7 ;
            rom[36286] = 8'h00 ;
            rom[36287] = 8'he7 ;
            rom[36288] = 8'hf8 ;
            rom[36289] = 8'h03 ;
            rom[36290] = 8'hfd ;
            rom[36291] = 8'he4 ;
            rom[36292] = 8'h01 ;
            rom[36293] = 8'h1f ;
            rom[36294] = 8'hd0 ;
            rom[36295] = 8'hff ;
            rom[36296] = 8'h15 ;
            rom[36297] = 8'h15 ;
            rom[36298] = 8'h05 ;
            rom[36299] = 8'hee ;
            rom[36300] = 8'he4 ;
            rom[36301] = 8'hee ;
            rom[36302] = 8'hee ;
            rom[36303] = 8'hf1 ;
            rom[36304] = 8'hf2 ;
            rom[36305] = 8'hcf ;
            rom[36306] = 8'h0d ;
            rom[36307] = 8'hd3 ;
            rom[36308] = 8'he4 ;
            rom[36309] = 8'hf8 ;
            rom[36310] = 8'hf1 ;
            rom[36311] = 8'hfd ;
            rom[36312] = 8'hf3 ;
            rom[36313] = 8'h0f ;
            rom[36314] = 8'hf7 ;
            rom[36315] = 8'hea ;
            rom[36316] = 8'h0c ;
            rom[36317] = 8'hf4 ;
            rom[36318] = 8'hac ;
            rom[36319] = 8'hbf ;
            rom[36320] = 8'hd1 ;
            rom[36321] = 8'hf8 ;
            rom[36322] = 8'h15 ;
            rom[36323] = 8'hee ;
            rom[36324] = 8'h03 ;
            rom[36325] = 8'heb ;
            rom[36326] = 8'h00 ;
            rom[36327] = 8'hf3 ;
            rom[36328] = 8'he2 ;
            rom[36329] = 8'h1a ;
            rom[36330] = 8'he3 ;
            rom[36331] = 8'hef ;
            rom[36332] = 8'he1 ;
            rom[36333] = 8'hf5 ;
            rom[36334] = 8'hf4 ;
            rom[36335] = 8'h11 ;
            rom[36336] = 8'hf4 ;
            rom[36337] = 8'h14 ;
            rom[36338] = 8'h12 ;
            rom[36339] = 8'hda ;
            rom[36340] = 8'h00 ;
            rom[36341] = 8'h0d ;
            rom[36342] = 8'hfe ;
            rom[36343] = 8'h04 ;
            rom[36344] = 8'he7 ;
            rom[36345] = 8'h00 ;
            rom[36346] = 8'hda ;
            rom[36347] = 8'h1a ;
            rom[36348] = 8'he9 ;
            rom[36349] = 8'h1b ;
            rom[36350] = 8'hf0 ;
            rom[36351] = 8'he9 ;
            rom[36352] = 8'h05 ;
            rom[36353] = 8'heb ;
            rom[36354] = 8'he9 ;
            rom[36355] = 8'hee ;
            rom[36356] = 8'hf0 ;
            rom[36357] = 8'h00 ;
            rom[36358] = 8'h20 ;
            rom[36359] = 8'hee ;
            rom[36360] = 8'he5 ;
            rom[36361] = 8'hc9 ;
            rom[36362] = 8'h10 ;
            rom[36363] = 8'heb ;
            rom[36364] = 8'hdd ;
            rom[36365] = 8'hf7 ;
            rom[36366] = 8'h09 ;
            rom[36367] = 8'h05 ;
            rom[36368] = 8'h09 ;
            rom[36369] = 8'h0b ;
            rom[36370] = 8'he3 ;
            rom[36371] = 8'hde ;
            rom[36372] = 8'he0 ;
            rom[36373] = 8'h04 ;
            rom[36374] = 8'h16 ;
            rom[36375] = 8'h01 ;
            rom[36376] = 8'hb6 ;
            rom[36377] = 8'ha3 ;
            rom[36378] = 8'h0f ;
            rom[36379] = 8'hf4 ;
            rom[36380] = 8'hf8 ;
            rom[36381] = 8'he8 ;
            rom[36382] = 8'hb3 ;
            rom[36383] = 8'hff ;
            rom[36384] = 8'hf1 ;
            rom[36385] = 8'h20 ;
            rom[36386] = 8'h18 ;
            rom[36387] = 8'hd7 ;
            rom[36388] = 8'hf8 ;
            rom[36389] = 8'h01 ;
            rom[36390] = 8'hf6 ;
            rom[36391] = 8'hf6 ;
            rom[36392] = 8'h1a ;
            rom[36393] = 8'hf3 ;
            rom[36394] = 8'hf5 ;
            rom[36395] = 8'hfc ;
            rom[36396] = 8'he4 ;
            rom[36397] = 8'hec ;
            rom[36398] = 8'hed ;
            rom[36399] = 8'h13 ;
            rom[36400] = 8'hfb ;
            rom[36401] = 8'hd3 ;
            rom[36402] = 8'hf5 ;
            rom[36403] = 8'h0b ;
            rom[36404] = 8'he8 ;
            rom[36405] = 8'he8 ;
            rom[36406] = 8'hfd ;
            rom[36407] = 8'hfa ;
            rom[36408] = 8'h0c ;
            rom[36409] = 8'hdb ;
            rom[36410] = 8'he8 ;
            rom[36411] = 8'hfb ;
            rom[36412] = 8'h01 ;
            rom[36413] = 8'hfc ;
            rom[36414] = 8'he6 ;
            rom[36415] = 8'h13 ;
            rom[36416] = 8'he1 ;
            rom[36417] = 8'hea ;
            rom[36418] = 8'hde ;
            rom[36419] = 8'hfd ;
            rom[36420] = 8'he2 ;
            rom[36421] = 8'hf5 ;
            rom[36422] = 8'he7 ;
            rom[36423] = 8'h14 ;
            rom[36424] = 8'h0c ;
            rom[36425] = 8'hf6 ;
            rom[36426] = 8'h07 ;
            rom[36427] = 8'h04 ;
            rom[36428] = 8'he7 ;
            rom[36429] = 8'h10 ;
            rom[36430] = 8'hff ;
            rom[36431] = 8'h17 ;
            rom[36432] = 8'h03 ;
            rom[36433] = 8'h0c ;
            rom[36434] = 8'hfe ;
            rom[36435] = 8'hfa ;
            rom[36436] = 8'h14 ;
            rom[36437] = 8'he4 ;
            rom[36438] = 8'h01 ;
            rom[36439] = 8'hf3 ;
            rom[36440] = 8'hea ;
            rom[36441] = 8'hf2 ;
            rom[36442] = 8'h10 ;
            rom[36443] = 8'h13 ;
            rom[36444] = 8'hd2 ;
            rom[36445] = 8'hf6 ;
            rom[36446] = 8'h0e ;
            rom[36447] = 8'hf8 ;
            rom[36448] = 8'h07 ;
            rom[36449] = 8'h1d ;
            rom[36450] = 8'h03 ;
            rom[36451] = 8'h06 ;
            rom[36452] = 8'he7 ;
            rom[36453] = 8'hc9 ;
            rom[36454] = 8'h10 ;
            rom[36455] = 8'hf7 ;
            rom[36456] = 8'h02 ;
            rom[36457] = 8'h16 ;
            rom[36458] = 8'hf9 ;
            rom[36459] = 8'h0d ;
            rom[36460] = 8'h03 ;
            rom[36461] = 8'hf7 ;
            rom[36462] = 8'h1c ;
            rom[36463] = 8'hfa ;
            rom[36464] = 8'h0f ;
            rom[36465] = 8'h07 ;
            rom[36466] = 8'h0f ;
            rom[36467] = 8'hfe ;
            rom[36468] = 8'hfe ;
            rom[36469] = 8'he7 ;
            rom[36470] = 8'hed ;
            rom[36471] = 8'h18 ;
            rom[36472] = 8'h1c ;
            rom[36473] = 8'hfb ;
            rom[36474] = 8'hd6 ;
            rom[36475] = 8'h15 ;
            rom[36476] = 8'hf1 ;
            rom[36477] = 8'h03 ;
            rom[36478] = 8'h0f ;
            rom[36479] = 8'hbf ;
            rom[36480] = 8'h07 ;
            rom[36481] = 8'hf4 ;
            rom[36482] = 8'hfd ;
            rom[36483] = 8'hfd ;
            rom[36484] = 8'h0a ;
            rom[36485] = 8'hed ;
            rom[36486] = 8'h2c ;
            rom[36487] = 8'hef ;
            rom[36488] = 8'h07 ;
            rom[36489] = 8'hf2 ;
            rom[36490] = 8'hf7 ;
            rom[36491] = 8'hec ;
            rom[36492] = 8'h01 ;
            rom[36493] = 8'hb1 ;
            rom[36494] = 8'h0b ;
            rom[36495] = 8'hef ;
            rom[36496] = 8'h0d ;
            rom[36497] = 8'hc5 ;
            rom[36498] = 8'hf7 ;
            rom[36499] = 8'h07 ;
            rom[36500] = 8'h04 ;
            rom[36501] = 8'hfd ;
            rom[36502] = 8'hf4 ;
            rom[36503] = 8'hf9 ;
            rom[36504] = 8'hef ;
            rom[36505] = 8'hfd ;
            rom[36506] = 8'hf9 ;
            rom[36507] = 8'hfa ;
            rom[36508] = 8'h00 ;
            rom[36509] = 8'h09 ;
            rom[36510] = 8'hf8 ;
            rom[36511] = 8'hf3 ;
            rom[36512] = 8'h09 ;
            rom[36513] = 8'h10 ;
            rom[36514] = 8'h03 ;
            rom[36515] = 8'he0 ;
            rom[36516] = 8'hc9 ;
            rom[36517] = 8'h06 ;
            rom[36518] = 8'h05 ;
            rom[36519] = 8'h18 ;
            rom[36520] = 8'hd9 ;
            rom[36521] = 8'hfd ;
            rom[36522] = 8'h21 ;
            rom[36523] = 8'h03 ;
            rom[36524] = 8'h08 ;
            rom[36525] = 8'h14 ;
            rom[36526] = 8'hf2 ;
            rom[36527] = 8'hf2 ;
            rom[36528] = 8'hec ;
            rom[36529] = 8'hfb ;
            rom[36530] = 8'h04 ;
            rom[36531] = 8'hae ;
            rom[36532] = 8'hbe ;
            rom[36533] = 8'h02 ;
            rom[36534] = 8'hea ;
            rom[36535] = 8'hdf ;
            rom[36536] = 8'hf6 ;
            rom[36537] = 8'h09 ;
            rom[36538] = 8'h0a ;
            rom[36539] = 8'hea ;
            rom[36540] = 8'h1a ;
            rom[36541] = 8'hf6 ;
            rom[36542] = 8'hf5 ;
            rom[36543] = 8'hbb ;
            rom[36544] = 8'hf0 ;
            rom[36545] = 8'hd5 ;
            rom[36546] = 8'hec ;
            rom[36547] = 8'hf7 ;
            rom[36548] = 8'he1 ;
            rom[36549] = 8'hf3 ;
            rom[36550] = 8'hce ;
            rom[36551] = 8'hf8 ;
            rom[36552] = 8'hf1 ;
            rom[36553] = 8'hed ;
            rom[36554] = 8'h19 ;
            rom[36555] = 8'hd7 ;
            rom[36556] = 8'hf9 ;
            rom[36557] = 8'he4 ;
            rom[36558] = 8'hf1 ;
            rom[36559] = 8'he9 ;
            rom[36560] = 8'hf8 ;
            rom[36561] = 8'he8 ;
            rom[36562] = 8'hf7 ;
            rom[36563] = 8'hdc ;
            rom[36564] = 8'h15 ;
            rom[36565] = 8'he2 ;
            rom[36566] = 8'h05 ;
            rom[36567] = 8'he1 ;
            rom[36568] = 8'h00 ;
            rom[36569] = 8'hf0 ;
            rom[36570] = 8'h29 ;
            rom[36571] = 8'h0c ;
            rom[36572] = 8'hfd ;
            rom[36573] = 8'he3 ;
            rom[36574] = 8'hce ;
            rom[36575] = 8'hef ;
            rom[36576] = 8'h0e ;
            rom[36577] = 8'hef ;
            rom[36578] = 8'hd5 ;
            rom[36579] = 8'hed ;
            rom[36580] = 8'h0e ;
            rom[36581] = 8'h09 ;
            rom[36582] = 8'hf5 ;
            rom[36583] = 8'hea ;
            rom[36584] = 8'h01 ;
            rom[36585] = 8'heb ;
            rom[36586] = 8'hc3 ;
            rom[36587] = 8'hfe ;
            rom[36588] = 8'h08 ;
            rom[36589] = 8'h0c ;
            rom[36590] = 8'h0f ;
            rom[36591] = 8'hf5 ;
            rom[36592] = 8'h06 ;
            rom[36593] = 8'hf7 ;
            rom[36594] = 8'hec ;
            rom[36595] = 8'h14 ;
            rom[36596] = 8'hcf ;
            rom[36597] = 8'h0b ;
            rom[36598] = 8'he1 ;
            rom[36599] = 8'h03 ;
            rom[36600] = 8'he8 ;
            rom[36601] = 8'hcc ;
            rom[36602] = 8'hee ;
            rom[36603] = 8'h02 ;
            rom[36604] = 8'haf ;
            rom[36605] = 8'hb2 ;
            rom[36606] = 8'h11 ;
            rom[36607] = 8'h0c ;
            rom[36608] = 8'h1c ;
            rom[36609] = 8'h0c ;
            rom[36610] = 8'h0a ;
            rom[36611] = 8'h03 ;
            rom[36612] = 8'he6 ;
            rom[36613] = 8'h0f ;
            rom[36614] = 8'h00 ;
            rom[36615] = 8'hf4 ;
            rom[36616] = 8'hfc ;
            rom[36617] = 8'hfc ;
            rom[36618] = 8'h07 ;
            rom[36619] = 8'he5 ;
            rom[36620] = 8'hfe ;
            rom[36621] = 8'hca ;
            rom[36622] = 8'h05 ;
            rom[36623] = 8'h02 ;
            rom[36624] = 8'h06 ;
            rom[36625] = 8'h05 ;
            rom[36626] = 8'hfa ;
            rom[36627] = 8'hdd ;
            rom[36628] = 8'h0f ;
            rom[36629] = 8'h0f ;
            rom[36630] = 8'h17 ;
            rom[36631] = 8'h01 ;
            rom[36632] = 8'hf2 ;
            rom[36633] = 8'h1d ;
            rom[36634] = 8'hf2 ;
            rom[36635] = 8'h01 ;
            rom[36636] = 8'hfa ;
            rom[36637] = 8'hfe ;
            rom[36638] = 8'h19 ;
            rom[36639] = 8'h14 ;
            rom[36640] = 8'hf2 ;
            rom[36641] = 8'hfa ;
            rom[36642] = 8'hf6 ;
            rom[36643] = 8'h17 ;
            rom[36644] = 8'h14 ;
            rom[36645] = 8'hef ;
            rom[36646] = 8'hf5 ;
            rom[36647] = 8'hf8 ;
            rom[36648] = 8'hea ;
            rom[36649] = 8'he4 ;
            rom[36650] = 8'he4 ;
            rom[36651] = 8'h10 ;
            rom[36652] = 8'h05 ;
            rom[36653] = 8'hf4 ;
            rom[36654] = 8'hde ;
            rom[36655] = 8'h01 ;
            rom[36656] = 8'he3 ;
            rom[36657] = 8'h04 ;
            rom[36658] = 8'h19 ;
            rom[36659] = 8'hd6 ;
            rom[36660] = 8'hf4 ;
            rom[36661] = 8'h06 ;
            rom[36662] = 8'hd2 ;
            rom[36663] = 8'h0d ;
            rom[36664] = 8'h0c ;
            rom[36665] = 8'h19 ;
            rom[36666] = 8'hfd ;
            rom[36667] = 8'heb ;
            rom[36668] = 8'h17 ;
            rom[36669] = 8'h05 ;
            rom[36670] = 8'h16 ;
            rom[36671] = 8'hf6 ;
            rom[36672] = 8'hd7 ;
            rom[36673] = 8'hed ;
            rom[36674] = 8'he1 ;
            rom[36675] = 8'hf3 ;
            rom[36676] = 8'h23 ;
            rom[36677] = 8'h23 ;
            rom[36678] = 8'hea ;
            rom[36679] = 8'h00 ;
            rom[36680] = 8'hf5 ;
            rom[36681] = 8'h0f ;
            rom[36682] = 8'h07 ;
            rom[36683] = 8'hf0 ;
            rom[36684] = 8'h0c ;
            rom[36685] = 8'hd4 ;
            rom[36686] = 8'hde ;
            rom[36687] = 8'hd6 ;
            rom[36688] = 8'h01 ;
            rom[36689] = 8'hd7 ;
            rom[36690] = 8'he9 ;
            rom[36691] = 8'hda ;
            rom[36692] = 8'hee ;
            rom[36693] = 8'h06 ;
            rom[36694] = 8'hed ;
            rom[36695] = 8'hff ;
            rom[36696] = 8'hf3 ;
            rom[36697] = 8'h17 ;
            rom[36698] = 8'h03 ;
            rom[36699] = 8'hc0 ;
            rom[36700] = 8'hf0 ;
            rom[36701] = 8'he9 ;
            rom[36702] = 8'h16 ;
            rom[36703] = 8'hfc ;
            rom[36704] = 8'he3 ;
            rom[36705] = 8'h00 ;
            rom[36706] = 8'hf8 ;
            rom[36707] = 8'hf3 ;
            rom[36708] = 8'hcf ;
            rom[36709] = 8'hf5 ;
            rom[36710] = 8'hed ;
            rom[36711] = 8'h05 ;
            rom[36712] = 8'h04 ;
            rom[36713] = 8'h17 ;
            rom[36714] = 8'hd4 ;
            rom[36715] = 8'hfe ;
            rom[36716] = 8'he9 ;
            rom[36717] = 8'h01 ;
            rom[36718] = 8'h05 ;
            rom[36719] = 8'hed ;
            rom[36720] = 8'he7 ;
            rom[36721] = 8'hfa ;
            rom[36722] = 8'hf1 ;
            rom[36723] = 8'hfb ;
            rom[36724] = 8'h19 ;
            rom[36725] = 8'he1 ;
            rom[36726] = 8'hff ;
            rom[36727] = 8'hf7 ;
            rom[36728] = 8'hc7 ;
            rom[36729] = 8'hcc ;
            rom[36730] = 8'he7 ;
            rom[36731] = 8'h25 ;
            rom[36732] = 8'he0 ;
            rom[36733] = 8'hfe ;
            rom[36734] = 8'h0d ;
            rom[36735] = 8'h10 ;
            rom[36736] = 8'hfe ;
            rom[36737] = 8'hc5 ;
            rom[36738] = 8'hf3 ;
            rom[36739] = 8'hee ;
            rom[36740] = 8'hec ;
            rom[36741] = 8'hf8 ;
            rom[36742] = 8'hf6 ;
            rom[36743] = 8'h22 ;
            rom[36744] = 8'h01 ;
            rom[36745] = 8'h07 ;
            rom[36746] = 8'h15 ;
            rom[36747] = 8'hca ;
            rom[36748] = 8'hf8 ;
            rom[36749] = 8'h2b ;
            rom[36750] = 8'h2b ;
            rom[36751] = 8'hb5 ;
            rom[36752] = 8'h06 ;
            rom[36753] = 8'h11 ;
            rom[36754] = 8'hfb ;
            rom[36755] = 8'h0b ;
            rom[36756] = 8'hcd ;
            rom[36757] = 8'he5 ;
            rom[36758] = 8'hed ;
            rom[36759] = 8'h01 ;
            rom[36760] = 8'h01 ;
            rom[36761] = 8'h06 ;
            rom[36762] = 8'h1b ;
            rom[36763] = 8'hf4 ;
            rom[36764] = 8'h08 ;
            rom[36765] = 8'h2c ;
            rom[36766] = 8'hd0 ;
            rom[36767] = 8'hea ;
            rom[36768] = 8'he5 ;
            rom[36769] = 8'hdf ;
            rom[36770] = 8'hef ;
            rom[36771] = 8'hd6 ;
            rom[36772] = 8'he2 ;
            rom[36773] = 8'hff ;
            rom[36774] = 8'h06 ;
            rom[36775] = 8'he7 ;
            rom[36776] = 8'hd5 ;
            rom[36777] = 8'hed ;
            rom[36778] = 8'he0 ;
            rom[36779] = 8'he2 ;
            rom[36780] = 8'hf5 ;
            rom[36781] = 8'h0b ;
            rom[36782] = 8'hdb ;
            rom[36783] = 8'heb ;
            rom[36784] = 8'h08 ;
            rom[36785] = 8'he4 ;
            rom[36786] = 8'h0d ;
            rom[36787] = 8'h14 ;
            rom[36788] = 8'hf0 ;
            rom[36789] = 8'he2 ;
            rom[36790] = 8'he3 ;
            rom[36791] = 8'hf6 ;
            rom[36792] = 8'hf3 ;
            rom[36793] = 8'hcf ;
            rom[36794] = 8'he9 ;
            rom[36795] = 8'h05 ;
            rom[36796] = 8'hab ;
            rom[36797] = 8'hfc ;
            rom[36798] = 8'hea ;
            rom[36799] = 8'hd9 ;
            rom[36800] = 8'h01 ;
            rom[36801] = 8'hf7 ;
            rom[36802] = 8'hf9 ;
            rom[36803] = 8'hea ;
            rom[36804] = 8'hfa ;
            rom[36805] = 8'hd2 ;
            rom[36806] = 8'hf9 ;
            rom[36807] = 8'hc9 ;
            rom[36808] = 8'h0a ;
            rom[36809] = 8'hbb ;
            rom[36810] = 8'h16 ;
            rom[36811] = 8'h12 ;
            rom[36812] = 8'hfc ;
            rom[36813] = 8'h03 ;
            rom[36814] = 8'hf6 ;
            rom[36815] = 8'h02 ;
            rom[36816] = 8'hf4 ;
            rom[36817] = 8'hf2 ;
            rom[36818] = 8'he0 ;
            rom[36819] = 8'hf0 ;
            rom[36820] = 8'hf6 ;
            rom[36821] = 8'h04 ;
            rom[36822] = 8'he2 ;
            rom[36823] = 8'h02 ;
            rom[36824] = 8'h0d ;
            rom[36825] = 8'hca ;
            rom[36826] = 8'hcd ;
            rom[36827] = 8'hfe ;
            rom[36828] = 8'h09 ;
            rom[36829] = 8'hef ;
            rom[36830] = 8'hfe ;
            rom[36831] = 8'h04 ;
            rom[36832] = 8'h07 ;
            rom[36833] = 8'hf0 ;
            rom[36834] = 8'he5 ;
            rom[36835] = 8'hfa ;
            rom[36836] = 8'he7 ;
            rom[36837] = 8'he4 ;
            rom[36838] = 8'hd2 ;
            rom[36839] = 8'h04 ;
            rom[36840] = 8'he0 ;
            rom[36841] = 8'h02 ;
            rom[36842] = 8'h26 ;
            rom[36843] = 8'h02 ;
            rom[36844] = 8'h0d ;
            rom[36845] = 8'hd8 ;
            rom[36846] = 8'hf3 ;
            rom[36847] = 8'h06 ;
            rom[36848] = 8'hdf ;
            rom[36849] = 8'hf5 ;
            rom[36850] = 8'hfa ;
            rom[36851] = 8'h1f ;
            rom[36852] = 8'hbc ;
            rom[36853] = 8'hf4 ;
            rom[36854] = 8'h06 ;
            rom[36855] = 8'h02 ;
            rom[36856] = 8'h05 ;
            rom[36857] = 8'h0d ;
            rom[36858] = 8'he9 ;
            rom[36859] = 8'hdf ;
            rom[36860] = 8'hd2 ;
            rom[36861] = 8'hf3 ;
            rom[36862] = 8'hd6 ;
            rom[36863] = 8'hea ;
        end
    always
        @(*)
        begin
            data = rom[addr] ;
        end
endmodule
